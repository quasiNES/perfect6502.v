module Perfect6502 ( 
    input  reset,
    input  ready,
    input  clock0,
    output clock1,
    output clock2,
    input irq,
    input nmi,
    input so,
    output sync,
    output readNotWrite,
    output [15:0] address,
    inout [7:0] data
);

    wire [1724:0] nodes;

    pull1 (nodes[0]);
    
    
    
    pull1 (nodes[3]);
    
    pull1 (nodes[4]);
    
    pull1 (nodes[5]);
    
    pull1 (nodes[6]);
    
    
    pull1 (nodes[8]);
    
    
    pull1 (nodes[10]);
    
    pull1 (nodes[11]);
    
    
    
    pull1 (nodes[14]);
    
    
    pull1 (nodes[16]);
    
    pull1 (nodes[17]);
    
    
    pull1 (nodes[19]);
    
    pull1 (nodes[20]);
    
    pull1 (nodes[21]);
    
    pull1 (nodes[22]);
    
    pull1 (nodes[23]);
    
    
    pull1 (nodes[25]);
    
    pull1 (nodes[26]);
    
    pull1 (nodes[27]);
    
    
    pull1 (nodes[29]);
    
    pull1 (nodes[30]);
    
    pull1 (nodes[31]);
    
    
    pull1 (nodes[33]);
    
    pull1 (nodes[34]);
    
    pull1 (nodes[35]);
    
    pull1 (nodes[36]);
    
    
    pull1 (nodes[38]);
    
    pull1 (nodes[39]);
    
    
    
    
    
    
    
    pull1 (nodes[46]);
    
    
    
    
    
    
    
    pull1 (nodes[53]);
    
    
    
    
    
    pull1 (nodes[58]);
    
    
    pull1 (nodes[60]);
    
    pull1 (nodes[61]);
    
    pull1 (nodes[62]);
    
    pull1 (nodes[63]);
    
    
    pull1 (nodes[65]);
    
    
    pull1 (nodes[67]);
    
    
    
    pull1 (nodes[70]);
    
    pull1 (nodes[71]);
    
    pull1 (nodes[72]);
    
    
    
    pull1 (nodes[75]);
    
    pull1 (nodes[76]);
    
    pull1 (nodes[77]);
    
    pull1 (nodes[78]);
    
    pull1 (nodes[79]);
    
    pull1 (nodes[80]);
    
    
    
    pull1 (nodes[83]);
    
    pull1 (nodes[84]);
    
    
    
    
    
    pull1 (nodes[89]);
    
    pull1 (nodes[90]);
    
    pull1 (nodes[91]);
    
    
    pull1 (nodes[93]);
    
    
    
    
    pull1 (nodes[97]);
    
    
    
    
    
    
    
    pull1 (nodes[104]);
    
    pull1 (nodes[105]);
    
    
    
    pull1 (nodes[108]);
    
    pull1 (nodes[109]);
    
    pull1 (nodes[110]);
    
    pull1 (nodes[111]);
    
    
    pull1 (nodes[113]);
    
    
    
    
    pull1 (nodes[117]);
    
    pull1 (nodes[118]);
    
    
    pull1 (nodes[120]);
    
    
    pull1 (nodes[122]);
    
    pull1 (nodes[123]);
    
    pull1 (nodes[124]);
    
    pull1 (nodes[125]);
    
    
    pull1 (nodes[127]);
    
    pull1 (nodes[128]);
    
    
    pull1 (nodes[130]);
    
    pull1 (nodes[131]);
    
    pull1 (nodes[132]);
    
    pull1 (nodes[133]);
    
    pull1 (nodes[134]);
    
    
    
    
    
    pull1 (nodes[139]);
    
    
    pull1 (nodes[141]);
    
    pull1 (nodes[142]);
    
    pull1 (nodes[143]);
    
    pull1 (nodes[144]);
    
    pull1 (nodes[145]);
    
    pull1 (nodes[146]);
    
    
    
    pull1 (nodes[149]);
    
    
    
    pull1 (nodes[152]);
    
    
    pull1 (nodes[154]);
    
    pull1 (nodes[155]);
    
    pull1 (nodes[156]);
    
    pull1 (nodes[157]);
    
    
    
    pull1 (nodes[160]);
    
    pull1 (nodes[161]);
    
    
    pull1 (nodes[163]);
    
    
    
    
    pull1 (nodes[167]);
    
    pull1 (nodes[168]);
    
    pull1 (nodes[169]);
    
    
    
    pull1 (nodes[172]);
    
    pull1 (nodes[173]);
    
    pull1 (nodes[174]);
    
    
    pull1 (nodes[176]);
    
    pull1 (nodes[177]);
    
    pull1 (nodes[178]);
    
    pull1 (nodes[179]);
    
    pull1 (nodes[180]);
    
    
    pull1 (nodes[182]);
    
    
    pull1 (nodes[184]);
    
    
    
    pull1 (nodes[187]);
    
    pull1 (nodes[188]);
    
    
    
    pull1 (nodes[191]);
    
    pull1 (nodes[192]);
    
    pull1 (nodes[193]);
    
    pull1 (nodes[194]);
    
    
    pull1 (nodes[196]);
    
    
    pull1 (nodes[198]);
    
    
    pull1 (nodes[200]);
    
    pull1 (nodes[201]);
    
    
    
    pull1 (nodes[204]);
    
    
    pull1 (nodes[206]);
    
    pull1 (nodes[207]);
    
    pull1 (nodes[208]);
    
    pull1 (nodes[209]);
    
    
    
    pull1 (nodes[212]);
    
    pull1 (nodes[213]);
    
    
    
    pull1 (nodes[216]);
    
    pull1 (nodes[217]);
    
    pull1 (nodes[218]);
    
    pull1 (nodes[219]);
    
    pull1 (nodes[220]);
    
    pull1 (nodes[221]);
    
    
    
    pull1 (nodes[224]);
    
    pull1 (nodes[225]);
    
    
    pull1 (nodes[227]);
    
    pull1 (nodes[228]);
    
    pull1 (nodes[229]);
    
    
    pull1 (nodes[231]);
    
    pull1 (nodes[232]);
    
    pull1 (nodes[233]);
    
    pull1 (nodes[234]);
    
    
    pull1 (nodes[236]);
    
    
    pull1 (nodes[238]);
    
    
    pull1 (nodes[240]);
    
    pull1 (nodes[241]);
    
    pull1 (nodes[242]);
    
    pull1 (nodes[243]);
    
    pull1 (nodes[244]);
    
    pull1 (nodes[245]);
    
    
    
    
    pull1 (nodes[249]);
    
    
    pull1 (nodes[251]);
    
    pull1 (nodes[252]);
    
    pull1 (nodes[253]);
    
    pull1 (nodes[254]);
    
    pull1 (nodes[255]);
    
    pull1 (nodes[256]);
    
    pull1 (nodes[257]);
    
    pull1 (nodes[258]);
    
    pull1 (nodes[259]);
    
    pull1 (nodes[260]);
    
    pull1 (nodes[261]);
    
    pull1 (nodes[262]);
    
    pull1 (nodes[263]);
    
    pull1 (nodes[264]);
    
    
    
    pull1 (nodes[267]);
    
    
    pull1 (nodes[269]);
    
    pull1 (nodes[270]);
    
    pull1 (nodes[271]);
    
    pull1 (nodes[272]);
    
    pull1 (nodes[273]);
    
    pull1 (nodes[274]);
    
    pull1 (nodes[275]);
    
    
    
    pull1 (nodes[278]);
    
    pull1 (nodes[279]);
    
    pull1 (nodes[280]);
    
    pull1 (nodes[281]);
    
    pull1 (nodes[282]);
    
    
    pull1 (nodes[284]);
    
    pull1 (nodes[285]);
    
    pull1 (nodes[286]);
    
    pull1 (nodes[287]);
    
    pull1 (nodes[288]);
    
    
    pull1 (nodes[290]);
    
    pull1 (nodes[291]);
    
    
    pull1 (nodes[293]);
    
    
    pull1 (nodes[295]);
    
    
    pull1 (nodes[297]);
    
    
    pull1 (nodes[299]);
    
    pull1 (nodes[300]);
    
    pull1 (nodes[301]);
    
    pull1 (nodes[302]);
    
    pull1 (nodes[303]);
    
    
    
    pull1 (nodes[306]);
    
    pull1 (nodes[307]);
    
    pull1 (nodes[308]);
    
    pull1 (nodes[309]);
    
    
    pull1 (nodes[311]);
    
    pull1 (nodes[312]);
    
    
    pull1 (nodes[314]);
    
    
    
    pull1 (nodes[317]);
    
    pull1 (nodes[318]);
    
    pull1 (nodes[319]);
    
    pull1 (nodes[320]);
    
    pull1 (nodes[321]);
    
    
    
    pull1 (nodes[324]);
    
    
    pull1 (nodes[326]);
    
    pull1 (nodes[327]);
    
    pull1 (nodes[328]);
    
    pull1 (nodes[329]);
    
    pull1 (nodes[330]);
    
    pull1 (nodes[331]);
    
    pull1 (nodes[332]);
    
    pull1 (nodes[333]);
    
    pull1 (nodes[334]);
    
    pull1 (nodes[335]);
    
    pull1 (nodes[336]);
    
    pull1 (nodes[337]);
    
    
    
    pull1 (nodes[340]);
    
    pull1 (nodes[341]);
    
    pull1 (nodes[342]);
    
    
    pull1 (nodes[344]);
    
    pull1 (nodes[345]);
    
    
    pull1 (nodes[347]);
    
    
    
    pull1 (nodes[350]);
    
    pull1 (nodes[351]);
    
    pull1 (nodes[352]);
    
    
    pull1 (nodes[354]);
    
    pull1 (nodes[355]);
    
    
    
    pull1 (nodes[358]);
    
    
    
    
    
    
    
    pull1 (nodes[365]);
    
    pull1 (nodes[366]);
    
    
    pull1 (nodes[368]);
    
    
    pull1 (nodes[370]);
    
    pull1 (nodes[371]);
    
    pull1 (nodes[372]);
    
    
    pull1 (nodes[374]);
    
    
    pull1 (nodes[376]);
    
    
    pull1 (nodes[378]);
    
    pull1 (nodes[379]);
    
    
    
    pull1 (nodes[382]);
    
    pull1 (nodes[383]);
    
    pull1 (nodes[384]);
    
    pull1 (nodes[385]);
    
    pull1 (nodes[386]);
    
    
    pull1 (nodes[388]);
    
    pull1 (nodes[389]);
    
    pull1 (nodes[390]);
    
    pull1 (nodes[391]);
    
    pull1 (nodes[392]);
    
    
    
    
    pull1 (nodes[396]);
    
    pull1 (nodes[397]);
    
    
    
    pull1 (nodes[400]);
    
    pull1 (nodes[401]);
    
    
    pull1 (nodes[403]);
    
    pull1 (nodes[404]);
    
    
    
    
    
    pull1 (nodes[409]);
    
    pull1 (nodes[410]);
    
    pull1 (nodes[411]);
    
    pull1 (nodes[412]);
    
    
    
    
    
    
    
    pull1 (nodes[419]);
    
    pull1 (nodes[420]);
    
    
    pull1 (nodes[422]);
    
    pull1 (nodes[423]);
    
    pull1 (nodes[424]);
    
    pull1 (nodes[425]);
    
    
    pull1 (nodes[427]);
    
    pull1 (nodes[428]);
    
    
    
    
    pull1 (nodes[432]);
    
    
    pull1 (nodes[434]);
    
    
    pull1 (nodes[436]);
    
    
    
    pull1 (nodes[439]);
    
    pull1 (nodes[440]);
    
    pull1 (nodes[441]);
    
    pull1 (nodes[442]);
    
    
    pull1 (nodes[444]);
    
    pull1 (nodes[445]);
    
    pull1 (nodes[446]);
    
    pull1 (nodes[447]);
    
    
    
    pull1 (nodes[450]);
    
    
    
    pull1 (nodes[453]);
    
    
    
    
    pull1 (nodes[457]);
    
    pull1 (nodes[458]);
    
    
    
    pull1 (nodes[461]);
    
    pull1 (nodes[462]);
    
    
    pull1 (nodes[464]);
    
    pull1 (nodes[465]);
    
    pull1 (nodes[466]);
    
    pull1 (nodes[467]);
    
    pull1 (nodes[468]);
    
    
    pull1 (nodes[470]);
    
    
    pull1 (nodes[472]);
    
    pull1 (nodes[473]);
    
    pull1 (nodes[474]);
    
    
    pull1 (nodes[476]);
    
    pull1 (nodes[477]);
    
    pull1 (nodes[478]);
    
    pull1 (nodes[479]);
    
    pull1 (nodes[480]);
    
    pull1 (nodes[481]);
    
    
    
    pull1 (nodes[484]);
    
    pull1 (nodes[485]);
    
    pull1 (nodes[486]);
    
    pull1 (nodes[487]);
    
    pull1 (nodes[488]);
    
    pull1 (nodes[489]);
    
    pull1 (nodes[490]);
    
    pull1 (nodes[491]);
    
    pull1 (nodes[492]);
    
    
    pull1 (nodes[494]);
    
    
    pull1 (nodes[496]);
    
    pull1 (nodes[497]);
    
    
    pull1 (nodes[499]);
    
    pull1 (nodes[500]);
    
    pull1 (nodes[501]);
    
    
    pull1 (nodes[503]);
    
    pull1 (nodes[504]);
    
    pull1 (nodes[505]);
    
    pull1 (nodes[506]);
    
    pull1 (nodes[507]);
    
    
    
    pull1 (nodes[510]);
    
    
    
    pull1 (nodes[513]);
    
    
    pull1 (nodes[515]);
    
    pull1 (nodes[516]);
    
    pull1 (nodes[517]);
    
    pull1 (nodes[518]);
    
    pull1 (nodes[519]);
    
    
    
    pull1 (nodes[522]);
    
    pull1 (nodes[523]);
    
    
    pull1 (nodes[525]);
    
    
    
    pull1 (nodes[528]);
    
    
    
    pull1 (nodes[531]);
    
    pull1 (nodes[532]);
    
    pull1 (nodes[533]);
    
    
    pull1 (nodes[535]);
    
    
    
    pull1 (nodes[538]);
    
    
    pull1 (nodes[540]);
    
    
    pull1 (nodes[542]);
    
    pull1 (nodes[543]);
    
    pull1 (nodes[544]);
    
    
    pull1 (nodes[546]);
    
    
    pull1 (nodes[548]);
    
    
    pull1 (nodes[550]);
    
    pull1 (nodes[551]);
    
    pull1 (nodes[552]);
    
    pull1 (nodes[553]);
    
    
    pull1 (nodes[555]);
    
    pull1 (nodes[556]);
    
    
    
    
    
    
    
    pull1 (nodes[563]);
    
    pull1 (nodes[564]);
    
    pull1 (nodes[565]);
    
    pull1 (nodes[566]);
    
    pull1 (nodes[567]);
    
    pull1 (nodes[568]);
    
    
    pull1 (nodes[570]);
    
    pull1 (nodes[571]);
    
    pull1 (nodes[572]);
    
    
    
    pull1 (nodes[575]);
    
    
    
    pull1 (nodes[578]);
    
    pull1 (nodes[579]);
    
    
    
    pull1 (nodes[582]);
    
    pull1 (nodes[583]);
    
    
    
    pull1 (nodes[586]);
    
    pull1 (nodes[587]);
    
    pull1 (nodes[588]);
    
    
    
    
    pull1 (nodes[592]);
    
    pull1 (nodes[593]);
    
    pull1 (nodes[594]);
    
    pull1 (nodes[595]);
    
    
    
    
    
    pull1 (nodes[600]);
    
    
    pull1 (nodes[602]);
    
    pull1 (nodes[603]);
    
    pull1 (nodes[604]);
    
    
    pull1 (nodes[606]);
    
    pull1 (nodes[607]);
    
    pull1 (nodes[608]);
    
    pull1 (nodes[609]);
    
    
    pull1 (nodes[611]);
    
    
    pull1 (nodes[613]);
    
    
    
    pull1 (nodes[616]);
    
    pull1 (nodes[617]);
    
    pull1 (nodes[618]);
    
    
    pull1 (nodes[620]);
    
    
    
    pull1 (nodes[623]);
    
    pull1 (nodes[624]);
    
    pull1 (nodes[625]);
    
    pull1 (nodes[626]);
    
    
    pull1 (nodes[628]);
    
    pull1 (nodes[629]);
    
    pull1 (nodes[630]);
    
    pull1 (nodes[631]);
    
    pull1 (nodes[632]);
    
    
    
    
    pull1 (nodes[636]);
    
    pull1 (nodes[637]);
    
    pull1 (nodes[638]);
    
    
    pull1 (nodes[640]);
    
    pull1 (nodes[641]);
    
    
    
    
    pull1 (nodes[645]);
    
    pull1 (nodes[646]);
    
    pull1 (nodes[647]);
    
    
    pull1 (nodes[649]);
    
    
    pull1 (nodes[651]);
    
    pull1 (nodes[652]);
    
    
    
    
    
    
    pull1 (nodes[658]);
    
    
    pull1 (nodes[660]);
    
    
    pull1 (nodes[662]);
    
    
    pull1 (nodes[664]);
    
    pull1 (nodes[665]);
    
    
    pull1 (nodes[667]);
    
    
    pull1 (nodes[669]);
    
    pull1 (nodes[670]);
    
    
    
    pull1 (nodes[673]);
    
    pull1 (nodes[674]);
    
    
    
    pull1 (nodes[677]);
    
    pull1 (nodes[678]);
    
    pull1 (nodes[679]);
    
    
    pull1 (nodes[681]);
    
    pull1 (nodes[682]);
    
    
    
    
    pull1 (nodes[686]);
    
    pull1 (nodes[687]);
    
    
    pull1 (nodes[689]);
    
    pull1 (nodes[690]);
    
    pull1 (nodes[691]);
    
    pull1 (nodes[692]);
    
    pull1 (nodes[693]);
    
    pull1 (nodes[694]);
    
    pull1 (nodes[695]);
    
    pull1 (nodes[696]);
    
    
    
    pull1 (nodes[699]);
    
    pull1 (nodes[700]);
    
    pull1 (nodes[701]);
    
    pull1 (nodes[702]);
    
    
    
    
    
    
    pull1 (nodes[708]);
    
    pull1 (nodes[709]);
    
    
    
    pull1 (nodes[712]);
    
    pull1 (nodes[713]);
    
    pull1 (nodes[714]);
    
    pull1 (nodes[715]);
    
    
    pull1 (nodes[717]);
    
    pull1 (nodes[718]);
    
    
    pull1 (nodes[720]);
    
    pull1 (nodes[721]);
    
    
    pull1 (nodes[723]);
    
    
    pull1 (nodes[725]);
    
    pull1 (nodes[726]);
    
    
    pull1 (nodes[728]);
    
    
    pull1 (nodes[730]);
    
    pull1 (nodes[731]);
    
    pull1 (nodes[732]);
    
    pull1 (nodes[733]);
    
    
    pull1 (nodes[735]);
    
    
    
    
    pull1 (nodes[739]);
    
    
    
    
    pull1 (nodes[743]);
    
    pull1 (nodes[744]);
    
    
    pull1 (nodes[746]);
    
    pull1 (nodes[747]);
    
    pull1 (nodes[748]);
    
    pull1 (nodes[749]);
    
    pull1 (nodes[750]);
    
    
    
    pull1 (nodes[753]);
    
    pull1 (nodes[754]);
    
    pull1 (nodes[755]);
    
    
    pull1 (nodes[757]);
    
    
    
    
    pull1 (nodes[761]);
    
    pull1 (nodes[762]);
    
    pull1 (nodes[763]);
    
    pull1 (nodes[764]);
    
    pull1 (nodes[765]);
    
    
    pull1 (nodes[767]);
    
    
    pull1 (nodes[769]);
    
    pull1 (nodes[770]);
    
    pull1 (nodes[771]);
    
    pull1 (nodes[772]);
    
    pull1 (nodes[773]);
    
    pull1 (nodes[774]);
    
    pull1 (nodes[775]);
    
    pull1 (nodes[776]);
    
    
    pull1 (nodes[778]);
    
    pull1 (nodes[779]);
    
    
    pull1 (nodes[781]);
    
    pull1 (nodes[782]);
    
    pull1 (nodes[783]);
    
    pull1 (nodes[784]);
    
    
    pull1 (nodes[786]);
    
    pull1 (nodes[787]);
    
    pull1 (nodes[788]);
    
    pull1 (nodes[789]);
    
    pull1 (nodes[790]);
    
    pull1 (nodes[791]);
    
    
    
    
    pull1 (nodes[795]);
    
    
    pull1 (nodes[797]);
    
    
    
    pull1 (nodes[800]);
    
    
    
    pull1 (nodes[803]);
    
    pull1 (nodes[804]);
    
    
    
    pull1 (nodes[807]);
    
    pull1 (nodes[808]);
    
    pull1 (nodes[809]);
    
    pull1 (nodes[810]);
    
    pull1 (nodes[811]);
    
    pull1 (nodes[812]);
    
    pull1 (nodes[813]);
    
    
    pull1 (nodes[815]);
    
    
    pull1 (nodes[817]);
    
    pull1 (nodes[818]);
    
    pull1 (nodes[819]);
    
    
    
    pull1 (nodes[822]);
    
    
    pull1 (nodes[824]);
    
    
    
    pull1 (nodes[827]);
    
    
    
    pull1 (nodes[830]);
    
    pull1 (nodes[831]);
    
    
    
    pull1 (nodes[834]);
    
    
    
    pull1 (nodes[837]);
    
    pull1 (nodes[838]);
    
    pull1 (nodes[839]);
    
    pull1 (nodes[840]);
    
    pull1 (nodes[841]);
    
    pull1 (nodes[842]);
    
    
    pull1 (nodes[844]);
    
    pull1 (nodes[845]);
    
    pull1 (nodes[846]);
    
    pull1 (nodes[847]);
    
    
    pull1 (nodes[849]);
    
    pull1 (nodes[850]);
    
    pull1 (nodes[851]);
    
    pull1 (nodes[852]);
    
    pull1 (nodes[853]);
    
    pull1 (nodes[854]);
    
    
    
    pull1 (nodes[857]);
    
    
    
    pull1 (nodes[860]);
    
    pull1 (nodes[861]);
    
    pull1 (nodes[862]);
    
    
    
    
    
    pull1 (nodes[867]);
    
    
    
    pull1 (nodes[870]);
    
    pull1 (nodes[871]);
    
    pull1 (nodes[872]);
    
    
    
    pull1 (nodes[875]);
    
    pull1 (nodes[876]);
    
    pull1 (nodes[877]);
    
    
    pull1 (nodes[879]);
    
    pull1 (nodes[880]);
    
    
    pull1 (nodes[882]);
    
    pull1 (nodes[883]);
    
    pull1 (nodes[884]);
    
    pull1 (nodes[885]);
    
    
    
    pull1 (nodes[888]);
    
    pull1 (nodes[889]);
    
    pull1 (nodes[890]);
    
    
    
    
    
    pull1 (nodes[895]);
    
    pull1 (nodes[896]);
    
    
    
    
    
    pull1 (nodes[901]);
    
    
    
    pull1 (nodes[904]);
    
    pull1 (nodes[905]);
    
    pull1 (nodes[906]);
    
    
    pull1 (nodes[908]);
    
    pull1 (nodes[909]);
    
    pull1 (nodes[910]);
    
    
    
    pull1 (nodes[913]);
    
    
    pull1 (nodes[915]);
    
    pull1 (nodes[916]);
    
    pull1 (nodes[917]);
    
    pull1 (nodes[918]);
    
    pull1 (nodes[919]);
    
    pull1 (nodes[920]);
    
    
    
    pull1 (nodes[923]);
    
    
    pull1 (nodes[925]);
    
    pull1 (nodes[926]);
    
    
    pull1 (nodes[928]);
    
    pull1 (nodes[929]);
    
    pull1 (nodes[930]);
    
    pull1 (nodes[931]);
    
    pull1 (nodes[932]);
    
    pull1 (nodes[933]);
    
    pull1 (nodes[934]);
    
    pull1 (nodes[935]);
    
    pull1 (nodes[936]);
    
    pull1 (nodes[937]);
    
    pull1 (nodes[938]);
    
    
    
    
    
    
    pull1 (nodes[944]);
    
    
    pull1 (nodes[946]);
    
    pull1 (nodes[947]);
    
    
    
    pull1 (nodes[950]);
    
    pull1 (nodes[951]);
    
    pull1 (nodes[952]);
    
    pull1 (nodes[953]);
    
    pull1 (nodes[954]);
    
    
    pull1 (nodes[956]);
    
    
    pull1 (nodes[958]);
    
    pull1 (nodes[959]);
    
    
    pull1 (nodes[961]);
    
    pull1 (nodes[962]);
    
    
    pull1 (nodes[964]);
    
    pull1 (nodes[965]);
    
    pull1 (nodes[966]);
    
    pull1 (nodes[967]);
    
    
    pull1 (nodes[969]);
    
    
    pull1 (nodes[971]);
    
    
    pull1 (nodes[973]);
    
    
    pull1 (nodes[975]);
    
    pull1 (nodes[976]);
    
    
    
    pull1 (nodes[979]);
    
    pull1 (nodes[980]);
    
    pull1 (nodes[981]);
    
    
    pull1 (nodes[983]);
    
    
    pull1 (nodes[985]);
    
    pull1 (nodes[986]);
    
    pull1 (nodes[987]);
    
    pull1 (nodes[988]);
    
    
    pull1 (nodes[990]);
    
    
    pull1 (nodes[992]);
    
    
    
    pull1 (nodes[995]);
    
    pull1 (nodes[996]);
    
    pull1 (nodes[997]);
    
    pull1 (nodes[998]);
    
    
    
    
    pull1 (nodes[1002]);
    
    pull1 (nodes[1003]);
    
    
    
    pull1 (nodes[1006]);
    
    pull1 (nodes[1007]);
    
    
    pull1 (nodes[1009]);
    
    pull1 (nodes[1010]);
    
    
    
    
    
    
    pull1 (nodes[1016]);
    
    pull1 (nodes[1017]);
    
    pull1 (nodes[1018]);
    
    pull1 (nodes[1019]);
    
    
    pull1 (nodes[1021]);
    
    
    pull1 (nodes[1023]);
    
    pull1 (nodes[1024]);
    
    pull1 (nodes[1025]);
    
    pull1 (nodes[1026]);
    
    
    pull1 (nodes[1028]);
    
    
    
    pull1 (nodes[1031]);
    
    pull1 (nodes[1032]);
    
    pull1 (nodes[1033]);
    
    pull1 (nodes[1034]);
    
    pull1 (nodes[1035]);
    
    
    pull1 (nodes[1037]);
    
    pull1 (nodes[1038]);
    
    pull1 (nodes[1039]);
    
    
    
    pull1 (nodes[1042]);
    
    pull1 (nodes[1043]);
    
    pull1 (nodes[1044]);
    
    pull1 (nodes[1045]);
    
    pull1 (nodes[1046]);
    
    pull1 (nodes[1047]);
    
    pull1 (nodes[1048]);
    
    
    pull1 (nodes[1050]);
    
    
    pull1 (nodes[1052]);
    
    
    pull1 (nodes[1054]);
    
    pull1 (nodes[1055]);
    
    pull1 (nodes[1056]);
    
    pull1 (nodes[1057]);
    
    
    
    
    
    
    pull1 (nodes[1063]);
    
    
    pull1 (nodes[1065]);
    
    pull1 (nodes[1066]);
    
    pull1 (nodes[1067]);
    
    
    pull1 (nodes[1069]);
    
    pull1 (nodes[1070]);
    
    
    
    pull1 (nodes[1073]);
    
    pull1 (nodes[1074]);
    
    pull1 (nodes[1075]);
    
    
    pull1 (nodes[1077]);
    
    
    pull1 (nodes[1079]);
    
    
    pull1 (nodes[1081]);
    
    pull1 (nodes[1082]);
    
    pull1 (nodes[1083]);
    
    pull1 (nodes[1084]);
    
    pull1 (nodes[1085]);
    
    pull1 (nodes[1086]);
    
    pull1 (nodes[1087]);
    
    pull1 (nodes[1088]);
    
    pull1 (nodes[1089]);
    
    pull1 (nodes[1090]);
    
    pull1 (nodes[1091]);
    
    
    pull1 (nodes[1093]);
    
    pull1 (nodes[1094]);
    
    
    pull1 (nodes[1096]);
    
    pull1 (nodes[1097]);
    
    
    pull1 (nodes[1099]);
    
    
    pull1 (nodes[1101]);
    
    
    
    
    
    pull1 (nodes[1106]);
    
    pull1 (nodes[1107]);
    
    
    pull1 (nodes[1109]);
    
    pull1 (nodes[1110]);
    
    pull1 (nodes[1111]);
    
    pull1 (nodes[1112]);
    
    
    pull1 (nodes[1114]);
    
    pull1 (nodes[1115]);
    
    pull1 (nodes[1116]);
    
    pull1 (nodes[1117]);
    
    
    pull1 (nodes[1119]);
    
    pull1 (nodes[1120]);
    
    
    pull1 (nodes[1122]);
    
    
    
    pull1 (nodes[1125]);
    
    
    pull1 (nodes[1127]);
    
    
    pull1 (nodes[1129]);
    
    pull1 (nodes[1130]);
    
    
    
    pull1 (nodes[1133]);
    
    pull1 (nodes[1134]);
    
    pull1 (nodes[1135]);
    
    
    pull1 (nodes[1137]);
    
    pull1 (nodes[1138]);
    
    
    
    pull1 (nodes[1141]);
    
    
    pull1 (nodes[1143]);
    
    pull1 (nodes[1144]);
    
    pull1 (nodes[1145]);
    
    pull1 (nodes[1146]);
    
    
    
    
    
    
    
    pull1 (nodes[1153]);
    
    pull1 (nodes[1154]);
    
    pull1 (nodes[1155]);
    
    
    pull1 (nodes[1157]);
    
    
    pull1 (nodes[1159]);
    
    
    
    
    
    pull1 (nodes[1164]);
    
    pull1 (nodes[1165]);
    
    pull1 (nodes[1166]);
    
    
    pull1 (nodes[1168]);
    
    pull1 (nodes[1169]);
    
    pull1 (nodes[1170]);
    
    
    
    pull1 (nodes[1173]);
    
    pull1 (nodes[1174]);
    
    pull1 (nodes[1175]);
    
    
    
    pull1 (nodes[1178]);
    
    pull1 (nodes[1179]);
    
    pull1 (nodes[1180]);
    
    pull1 (nodes[1181]);
    
    pull1 (nodes[1182]);
    
    
    pull1 (nodes[1184]);
    
    pull1 (nodes[1185]);
    
    
    pull1 (nodes[1187]);
    
    
    
    pull1 (nodes[1190]);
    
    
    pull1 (nodes[1192]);
    
    pull1 (nodes[1193]);
    
    pull1 (nodes[1194]);
    
    pull1 (nodes[1195]);
    
    pull1 (nodes[1196]);
    
    pull1 (nodes[1197]);
    
    
    pull1 (nodes[1199]);
    
    pull1 (nodes[1200]);
    
    
    pull1 (nodes[1202]);
    
    
    pull1 (nodes[1204]);
    
    pull1 (nodes[1205]);
    
    pull1 (nodes[1206]);
    
    pull1 (nodes[1207]);
    
    pull1 (nodes[1208]);
    
    pull1 (nodes[1209]);
    
    pull1 (nodes[1210]);
    
    pull1 (nodes[1211]);
    
    
    pull1 (nodes[1213]);
    
    pull1 (nodes[1214]);
    
    pull1 (nodes[1215]);
    
    
    pull1 (nodes[1217]);
    
    pull1 (nodes[1218]);
    
    pull1 (nodes[1219]);
    
    pull1 (nodes[1220]);
    
    
    pull1 (nodes[1222]);
    
    pull1 (nodes[1223]);
    
    pull1 (nodes[1224]);
    
    pull1 (nodes[1225]);
    
    pull1 (nodes[1226]);
    
    pull1 (nodes[1227]);
    
    pull1 (nodes[1228]);
    
    pull1 (nodes[1229]);
    
    pull1 (nodes[1230]);
    
    pull1 (nodes[1231]);
    
    pull1 (nodes[1232]);
    
    pull1 (nodes[1233]);
    
    
    
    pull1 (nodes[1236]);
    
    
    pull1 (nodes[1238]);
    
    pull1 (nodes[1239]);
    
    pull1 (nodes[1240]);
    
    pull1 (nodes[1241]);
    
    
    pull1 (nodes[1243]);
    
    pull1 (nodes[1244]);
    
    pull1 (nodes[1245]);
    
    pull1 (nodes[1246]);
    
    
    
    
    pull1 (nodes[1250]);
    
    pull1 (nodes[1251]);
    
    
    pull1 (nodes[1253]);
    
    
    pull1 (nodes[1255]);
    
    pull1 (nodes[1256]);
    
    pull1 (nodes[1257]);
    
    pull1 (nodes[1258]);
    
    pull1 (nodes[1259]);
    
    pull1 (nodes[1260]);
    
    pull1 (nodes[1261]);
    
    pull1 (nodes[1262]);
    
    
    
    pull1 (nodes[1265]);
    
    
    pull1 (nodes[1267]);
    
    pull1 (nodes[1268]);
    
    
    pull1 (nodes[1270]);
    
    pull1 (nodes[1271]);
    
    
    pull1 (nodes[1273]);
    
    
    pull1 (nodes[1275]);
    
    
    pull1 (nodes[1277]);
    
    
    
    
    pull1 (nodes[1281]);
    
    
    
    
    pull1 (nodes[1285]);
    
    pull1 (nodes[1286]);
    
    
    
    pull1 (nodes[1289]);
    
    pull1 (nodes[1290]);
    
    
    pull1 (nodes[1292]);
    
    pull1 (nodes[1293]);
    
    pull1 (nodes[1294]);
    
    pull1 (nodes[1295]);
    
    
    
    
    
    
    pull1 (nodes[1301]);
    
    
    pull1 (nodes[1303]);
    
    pull1 (nodes[1304]);
    
    pull1 (nodes[1305]);
    
    pull1 (nodes[1306]);
    
    
    pull1 (nodes[1308]);
    
    pull1 (nodes[1309]);
    
    
    pull1 (nodes[1311]);
    
    pull1 (nodes[1312]);
    
    pull1 (nodes[1313]);
    
    pull1 (nodes[1314]);
    
    pull1 (nodes[1315]);
    
    pull1 (nodes[1316]);
    
    pull1 (nodes[1317]);
    
    pull1 (nodes[1318]);
    
    pull1 (nodes[1319]);
    
    pull1 (nodes[1320]);
    
    
    
    pull1 (nodes[1323]);
    
    pull1 (nodes[1324]);
    
    
    
    pull1 (nodes[1327]);
    
    pull1 (nodes[1328]);
    
    pull1 (nodes[1329]);
    
    
    
    
    
    pull1 (nodes[1334]);
    
    pull1 (nodes[1335]);
    
    
    pull1 (nodes[1337]);
    
    
    pull1 (nodes[1339]);
    
    
    
    pull1 (nodes[1342]);
    
    pull1 (nodes[1343]);
    
    pull1 (nodes[1344]);
    
    pull1 (nodes[1345]);
    
    pull1 (nodes[1346]);
    
    pull1 (nodes[1347]);
    
    
    
    pull1 (nodes[1350]);
    
    
    pull1 (nodes[1352]);
    
    
    
    pull1 (nodes[1355]);
    
    pull1 (nodes[1356]);
    
    pull1 (nodes[1357]);
    
    pull1 (nodes[1358]);
    
    
    
    pull1 (nodes[1361]);
    
    
    pull1 (nodes[1363]);
    
    pull1 (nodes[1364]);
    
    
    
    
    pull1 (nodes[1368]);
    
    pull1 (nodes[1369]);
    
    pull1 (nodes[1370]);
    
    pull1 (nodes[1371]);
    
    pull1 (nodes[1372]);
    
    
    pull1 (nodes[1374]);
    
    pull1 (nodes[1375]);
    
    pull1 (nodes[1376]);
    
    pull1 (nodes[1377]);
    
    
    pull1 (nodes[1379]);
    
    pull1 (nodes[1380]);
    
    pull1 (nodes[1381]);
    
    pull1 (nodes[1382]);
    
    pull1 (nodes[1383]);
    
    pull1 (nodes[1384]);
    
    pull1 (nodes[1385]);
    
    pull1 (nodes[1386]);
    
    
    
    pull1 (nodes[1389]);
    
    
    pull1 (nodes[1391]);
    
    pull1 (nodes[1392]);
    
    
    pull1 (nodes[1394]);
    
    
    pull1 (nodes[1396]);
    
    
    pull1 (nodes[1398]);
    
    pull1 (nodes[1399]);
    
    pull1 (nodes[1400]);
    
    pull1 (nodes[1401]);
    
    pull1 (nodes[1402]);
    
    
    
    
    
    
    pull1 (nodes[1408]);
    
    
    pull1 (nodes[1410]);
    
    
    pull1 (nodes[1412]);
    
    pull1 (nodes[1413]);
    
    pull1 (nodes[1414]);
    
    pull1 (nodes[1415]);
    
    pull1 (nodes[1416]);
    
    
    
    pull1 (nodes[1419]);
    
    pull1 (nodes[1420]);
    
    pull1 (nodes[1421]);
    
    
    pull1 (nodes[1423]);
    
    
    pull1 (nodes[1425]);
    
    
    pull1 (nodes[1427]);
    
    pull1 (nodes[1428]);
    
    pull1 (nodes[1429]);
    
    pull1 (nodes[1430]);
    
    
    
    pull1 (nodes[1433]);
    
    pull1 (nodes[1434]);
    
    
    
    
    
    pull1 (nodes[1439]);
    
    pull1 (nodes[1440]);
    
    pull1 (nodes[1441]);
    
    
    
    pull1 (nodes[1444]);
    
    
    pull1 (nodes[1446]);
    
    
    pull1 (nodes[1448]);
    
    pull1 (nodes[1449]);
    
    
    
    
    pull1 (nodes[1453]);
    
    
    pull1 (nodes[1455]);
    
    
    pull1 (nodes[1457]);
    
    pull1 (nodes[1458]);
    
    pull1 (nodes[1459]);
    
    pull1 (nodes[1460]);
    
    pull1 (nodes[1461]);
    
    pull1 (nodes[1462]);
    
    pull1 (nodes[1463]);
    
    pull1 (nodes[1464]);
    
    pull1 (nodes[1465]);
    
    pull1 (nodes[1466]);
    
    
    
    pull1 (nodes[1469]);
    
    
    pull1 (nodes[1471]);
    
    
    
    pull1 (nodes[1474]);
    
    pull1 (nodes[1475]);
    
    pull1 (nodes[1476]);
    
    
    pull1 (nodes[1478]);
    
    
    
    pull1 (nodes[1481]);
    
    pull1 (nodes[1482]);
    
    
    pull1 (nodes[1484]);
    
    
    pull1 (nodes[1486]);
    
    pull1 (nodes[1487]);
    
    pull1 (nodes[1488]);
    
    
    
    pull1 (nodes[1491]);
    
    pull1 (nodes[1492]);
    
    
    pull1 (nodes[1494]);
    
    pull1 (nodes[1495]);
    
    pull1 (nodes[1496]);
    
    pull1 (nodes[1497]);
    
    
    pull1 (nodes[1499]);
    
    pull1 (nodes[1500]);
    
    
    pull1 (nodes[1502]);
    
    
    pull1 (nodes[1504]);
    
    
    pull1 (nodes[1506]);
    
    pull1 (nodes[1507]);
    
    
    
    
    pull1 (nodes[1511]);
    
    pull1 (nodes[1512]);
    
    
    
    
    
    pull1 (nodes[1517]);
    
    pull1 (nodes[1518]);
    
    pull1 (nodes[1519]);
    
    pull1 (nodes[1520]);
    
    pull1 (nodes[1521]);
    
    
    pull1 (nodes[1523]);
    
    pull1 (nodes[1524]);
    
    pull1 (nodes[1525]);
    
    pull1 (nodes[1526]);
    
    
    
    
    
    pull1 (nodes[1531]);
    
    
    
    pull1 (nodes[1534]);
    
    
    
    
    
    
    pull1 (nodes[1540]);
    
    pull1 (nodes[1541]);
    
    pull1 (nodes[1542]);
    
    pull1 (nodes[1543]);
    
    pull1 (nodes[1544]);
    
    
    
    
    pull1 (nodes[1548]);
    
    pull1 (nodes[1549]);
    
    
    
    pull1 (nodes[1552]);
    
    
    
    
    
    pull1 (nodes[1557]);
    
    
    
    pull1 (nodes[1560]);
    
    pull1 (nodes[1561]);
    
    pull1 (nodes[1562]);
    
    
    
    
    pull1 (nodes[1566]);
    
    pull1 (nodes[1567]);
    
    
    pull1 (nodes[1569]);
    
    
    pull1 (nodes[1571]);
    
    
    pull1 (nodes[1573]);
    
    
    pull1 (nodes[1575]);
    
    pull1 (nodes[1576]);
    
    
    pull1 (nodes[1578]);
    
    
    pull1 (nodes[1580]);
    
    
    pull1 (nodes[1582]);
    
    
    
    pull1 (nodes[1585]);
    
    pull1 (nodes[1586]);
    
    pull1 (nodes[1587]);
    
    pull1 (nodes[1588]);
    
    pull1 (nodes[1589]);
    
    
    
    pull1 (nodes[1592]);
    
    pull1 (nodes[1593]);
    
    pull1 (nodes[1594]);
    
    pull1 (nodes[1595]);
    
    pull1 (nodes[1596]);
    
    pull1 (nodes[1597]);
    
    
    pull1 (nodes[1599]);
    
    pull1 (nodes[1600]);
    
    pull1 (nodes[1601]);
    
    
    
    
    pull1 (nodes[1605]);
    
    
    
    
    
    pull1 (nodes[1610]);
    
    
    pull1 (nodes[1612]);
    
    pull1 (nodes[1613]);
    
    pull1 (nodes[1614]);
    
    
    
    
    pull1 (nodes[1618]);
    
    pull1 (nodes[1619]);
    
    
    pull1 (nodes[1621]);
    
    pull1 (nodes[1622]);
    
    pull1 (nodes[1623]);
    
    
    
    pull1 (nodes[1626]);
    
    
    pull1 (nodes[1628]);
    
    pull1 (nodes[1629]);
    
    
    pull1 (nodes[1631]);
    
    pull1 (nodes[1632]);
    
    
    pull1 (nodes[1634]);
    
    pull1 (nodes[1635]);
    
    
    pull1 (nodes[1637]);
    
    pull1 (nodes[1638]);
    
    
    pull1 (nodes[1640]);
    
    pull1 (nodes[1641]);
    
    pull1 (nodes[1642]);
    
    pull1 (nodes[1643]);
    
    
    
    pull1 (nodes[1646]);
    
    pull1 (nodes[1647]);
    
    
    pull1 (nodes[1649]);
    
    pull1 (nodes[1650]);
    
    
    
    
    pull1 (nodes[1654]);
    
    pull1 (nodes[1655]);
    
    
    pull1 (nodes[1657]);
    
    pull1 (nodes[1658]);
    
    
    pull1 (nodes[1660]);
    
    
    pull1 (nodes[1662]);
    
    pull1 (nodes[1663]);
    
    pull1 (nodes[1664]);
    
    pull1 (nodes[1665]);
    
    
    
    pull1 (nodes[1668]);
    
    
    
    pull1 (nodes[1671]);
    
    pull1 (nodes[1672]);
    
    
    
    
    pull1 (nodes[1676]);
    
    pull1 (nodes[1677]);
    
    
    
    
    
    pull1 (nodes[1682]);
    
    
    pull1 (nodes[1684]);
    
    
    
    pull1 (nodes[1687]);
    
    pull1 (nodes[1688]);
    
    pull1 (nodes[1689]);
    
    
    pull1 (nodes[1691]);
    
    
    
    pull1 (nodes[1694]);
    
    
    
    pull1 (nodes[1697]);
    
    
    
    
    pull1 (nodes[1701]);
    
    
    
    pull1 (nodes[1704]);
    
    pull1 (nodes[1705]);
    
    
    
    pull1 (nodes[1708]);
    
    pull1 (nodes[1709]);
    
    pull1 (nodes[1710]);
    
    pull1 (nodes[1711]);
    
    pull1 (nodes[1712]);
    
    
    pull1 (nodes[1714]);
    
    pull1 (nodes[1715]);
    
    pull1 (nodes[1716]);
    
    pull1 (nodes[1717]);
    
    pull1 (nodes[1718]);
    
    pull1 (nodes[1719]);
    
    pull1 (nodes[1720]);
    
    pull1 (nodes[1721]);
    
    pull1 (nodes[1722]);
    
    
    pull1 (nodes[1724]);
    
    

    tranif1 (nodes[217], nodes[558],  nodes[357]);
    tranif1 (nodes[349], nodes[657],  nodes[1608]);
    tranif1 (nodes[1146], nodes[558],  nodes[412]);
    tranif1 (nodes[943], nodes[558],  nodes[558]);
    tranif1 (nodes[657], nodes[230],  nodes[826]);
    tranif1 (nodes[1319], nodes[558],  nodes[82]);
    tranif1 (nodes[1514], nodes[289],  nodes[821]);
    tranif1 (nodes[1171], nodes[558],  nodes[558]);
    tranif1 (nodes[1199], nodes[558],  nodes[945]);
    tranif1 (nodes[1548], nodes[524],  nodes[710]);
    tranif1 (nodes[220], nodes[558],  nodes[190]);
    tranif1 (nodes[657], nodes[1247],  nodes[38]);
    tranif1 (nodes[558], nodes[189],  nodes[1248]);
    tranif1 (nodes[155], nodes[558],  nodes[1248]);
    tranif1 (nodes[346], nodes[558],  nodes[943]);
    tranif1 (nodes[657], nodes[148],  nodes[1140]);
    tranif1 (nodes[558], nodes[508],  nodes[1540]);
    tranif1 (nodes[1082], nodes[32],  nodes[710]);
    tranif1 (nodes[212], nodes[1451],  nodes[710]);
    tranif1 (nodes[534], nodes[558],  nodes[1247]);
    tranif1 (nodes[272], nodes[1162],  nodes[943]);
    tranif1 (nodes[418], nodes[983],  nodes[943]);
    tranif1 (nodes[468], nodes[1615],  nodes[248]);
    tranif1 (nodes[395], nodes[472],  nodes[248]);
    tranif1 (nodes[348], nodes[1495],  nodes[710]);
    tranif1 (nodes[558], nodes[1100],  nodes[1096]);
    tranif1 (nodes[1660], nodes[558],  nodes[1096]);
    tranif1 (nodes[657], nodes[855],  nodes[1096]);
    tranif1 (nodes[744], nodes[558],  nodes[1503]);
    tranif1 (nodes[558], nodes[1616],  nodes[44]);
    tranif1 (nodes[375], nodes[651],  nodes[78]);
    tranif1 (nodes[65], nodes[558],  nodes[78]);
    tranif1 (nodes[1378], nodes[928],  nodes[710]);
    tranif1 (nodes[74], nodes[1309],  nodes[710]);
    tranif1 (nodes[115], nodes[518],  nodes[943]);
    tranif1 (nodes[31], nodes[558],  nodes[32]);
    tranif1 (nodes[657], nodes[1405],  nodes[943]);
    tranif1 (nodes[1603], nodes[973],  nodes[943]);
    tranif1 (nodes[558], nodes[510],  nodes[347]);
    tranif1 (nodes[883], nodes[1667],  nodes[710]);
    tranif1 (nodes[558], nodes[1456],  nodes[706]);
    tranif1 (nodes[558], nodes[307],  nodes[1174]);
    tranif1 (nodes[409], nodes[558],  nodes[1622]);
    tranif1 (nodes[558], nodes[25],  nodes[192]);
    tranif1 (nodes[606], nodes[558],  nodes[1490]);
    tranif1 (nodes[767], nodes[1148],  nodes[943]);
    tranif1 (nodes[1248], nodes[1150],  nodes[549]);
    tranif1 (nodes[1332], nodes[1287],  nodes[549]);
    tranif1 (nodes[1188], nodes[1680],  nodes[549]);
    tranif1 (nodes[1405], nodes[1142],  nodes[549]);
    tranif1 (nodes[558], nodes[794],  nodes[353]);
    tranif1 (nodes[558], nodes[794],  nodes[353]);
    tranif1 (nodes[1700], nodes[558],  nodes[593]);
    tranif1 (nodes[54], nodes[1167],  nodes[549]);
    tranif1 (nodes[1362], nodes[613],  nodes[600]);
    tranif1 (nodes[166], nodes[530],  nodes[549]);
    tranif1 (nodes[1336], nodes[1627],  nodes[549]);
    tranif1 (nodes[1400], nodes[558],  nodes[948]);
    tranif1 (nodes[480], nodes[1092],  nodes[264]);
    tranif1 (nodes[558], nodes[632],  nodes[1582]);
    tranif1 (nodes[923], nodes[558],  nodes[584]);
    tranif1 (nodes[136], nodes[274],  nodes[1003]);
    tranif1 (nodes[558], nodes[860],  nodes[1003]);
    tranif1 (nodes[1527], nodes[1347],  nodes[943]);
    tranif1 (nodes[331], nodes[558],  nodes[68]);
    tranif1 (nodes[558], nodes[945],  nodes[558]);
    tranif1 (nodes[1495], nodes[1644],  nodes[1457]);
    tranif1 (nodes[558], nodes[1066],  nodes[1485]);
    tranif1 (nodes[1066], nodes[558],  nodes[1485]);
    tranif1 (nodes[558], nodes[1066],  nodes[1485]);
    tranif1 (nodes[1622], nodes[558],  nodes[1077]);
    tranif1 (nodes[558], nodes[667],  nodes[1077]);
    tranif1 (nodes[1336], nodes[115],  nodes[325]);
    tranif1 (nodes[785], nodes[920],  nodes[710]);
    tranif1 (nodes[558], nodes[748],  nodes[1318]);
    tranif1 (nodes[657], nodes[304],  nodes[362]);
    tranif1 (nodes[657], nodes[421],  nodes[127]);
    tranif1 (nodes[1405], nodes[989],  nodes[325]);
    tranif1 (nodes[790], nodes[558],  nodes[53]);
    tranif1 (nodes[1068], nodes[558],  nodes[763]);
    tranif1 (nodes[147], nodes[558],  nodes[1088]);
    tranif1 (nodes[1463], nodes[558],  nodes[1088]);
    tranif1 (nodes[493], nodes[1370],  nodes[1042]);
    tranif1 (nodes[1421], nodes[1473],  nodes[1042]);
    tranif1 (nodes[443], nodes[513],  nodes[943]);
    tranif1 (nodes[1646], nodes[1673],  nodes[943]);
    tranif1 (nodes[1516], nodes[490],  nodes[943]);
    tranif1 (nodes[558], nodes[856],  nodes[311]);
    tranif1 (nodes[558], nodes[835],  nodes[311]);
    tranif1 (nodes[1158], nodes[558],  nodes[783]);
    tranif1 (nodes[1704], nodes[558],  nodes[783]);
    tranif1 (nodes[1253], nodes[558],  nodes[783]);
    tranif1 (nodes[558], nodes[230],  nodes[381]);
    tranif1 (nodes[558], nodes[230],  nodes[381]);
    tranif1 (nodes[558], nodes[230],  nodes[381]);
    tranif1 (nodes[230], nodes[558],  nodes[381]);
    tranif1 (nodes[558], nodes[230],  nodes[381]);
    tranif1 (nodes[230], nodes[558],  nodes[381]);
    tranif1 (nodes[558], nodes[230],  nodes[381]);
    tranif1 (nodes[1343], nodes[558],  nodes[152]);
    tranif1 (nodes[558], nodes[371],  nodes[555]);
    tranif1 (nodes[207], nodes[558],  nodes[810]);
    tranif1 (nodes[558], nodes[501],  nodes[819]);
    tranif1 (nodes[558], nodes[1138],  nodes[1148]);
    tranif1 (nodes[672], nodes[657],  nodes[963]);
    tranif1 (nodes[558], nodes[202],  nodes[967]);
    tranif1 (nodes[558], nodes[972],  nodes[1691]);
    tranif1 (nodes[558], nodes[1563],  nodes[1342]);
    tranif1 (nodes[558], nodes[844],  nodes[786]);
    tranif1 (nodes[1296], nodes[657],  nodes[422]);
    tranif1 (nodes[558], nodes[1346],  nodes[422]);
    tranif1 (nodes[558], nodes[359],  nodes[422]);
    tranif1 (nodes[558], nodes[1680],  nodes[984]);
    tranif1 (nodes[365], nodes[558],  nodes[1410]);
    tranif1 (nodes[1145], nodes[558],  nodes[403]);
    tranif1 (nodes[558], nodes[746],  nodes[527]);
    tranif1 (nodes[1372], nodes[972],  nodes[1610]);
    tranif1 (nodes[1497], nodes[653],  nodes[710]);
    tranif1 (nodes[558], nodes[489],  nodes[429]);
    tranif1 (nodes[10], nodes[558],  nodes[467]);
    tranif1 (nodes[558], nodes[692],  nodes[460]);
    tranif1 (nodes[1647], nodes[558],  nodes[536]);
    tranif1 (nodes[558], nodes[1358],  nodes[917]);
    tranif1 (nodes[514], nodes[429],  nodes[821]);
    tranif1 (nodes[1268], nodes[558],  nodes[744]);
    tranif1 (nodes[1570], nodes[430],  nodes[710]);
    tranif1 (nodes[393], nodes[1179],  nodes[943]);
    tranif1 (nodes[1188], nodes[998],  nodes[1700]);
    tranif1 (nodes[1287], nodes[1389],  nodes[1700]);
    tranif1 (nodes[1462], nodes[558],  nodes[1369]);
    tranif1 (nodes[438], nodes[657],  nodes[1369]);
    tranif1 (nodes[816], nodes[558],  nodes[925]);
    tranif1 (nodes[1001], nodes[721],  nodes[1700]);
    tranif1 (nodes[1336], nodes[618],  nodes[1700]);
    tranif1 (nodes[558], nodes[1043],  nodes[818]);
    tranif1 (nodes[414], nodes[657],  nodes[818]);
    tranif1 (nodes[1405], nodes[3],  nodes[1700]);
    tranif1 (nodes[558], nodes[1426],  nodes[270]);
    tranif1 (nodes[1559], nodes[477],  nodes[1678]);
    tranif1 (nodes[1632], nodes[558],  nodes[1678]);
    tranif1 (nodes[1083], nodes[1590],  nodes[710]);
    tranif1 (nodes[1017], nodes[558],  nodes[589]);
    tranif1 (nodes[1066], nodes[1424],  nodes[710]);
    tranif1 (nodes[558], nodes[1455],  nodes[1420]);
    tranif1 (nodes[558], nodes[397],  nodes[1420]);
    tranif1 (nodes[558], nodes[789],  nodes[493]);
    tranif1 (nodes[558], nodes[884],  nodes[640]);
    tranif1 (nodes[624], nodes[558],  nodes[1108]);
    tranif1 (nodes[75], nodes[558],  nodes[154]);
    tranif1 (nodes[129], nodes[657],  nodes[154]);
    tranif1 (nodes[605], nodes[558],  nodes[787]);
    tranif1 (nodes[325], nodes[558],  nodes[1247]);
    tranif1 (nodes[558], nodes[604],  nodes[1582]);
    tranif1 (nodes[558], nodes[1010],  nodes[1670]);
    tranif1 (nodes[657], nodes[82],  nodes[798]);
    tranif1 (nodes[657], nodes[82],  nodes[798]);
    tranif1 (nodes[558], nodes[1264],  nodes[453]);
    tranif1 (nodes[558], nodes[567],  nodes[28]);
    tranif1 (nodes[1548], nodes[558],  nodes[121]);
    tranif1 (nodes[558], nodes[1225],  nodes[285]);
    tranif1 (nodes[70], nodes[558],  nodes[1134]);
    tranif1 (nodes[558], nodes[1366],  nodes[706]);
    tranif1 (nodes[558], nodes[952],  nodes[272]);
    tranif1 (nodes[558], nodes[426],  nodes[715]);
    tranif1 (nodes[558], nodes[914],  nodes[715]);
    tranif1 (nodes[739], nodes[711],  nodes[761]);
    tranif1 (nodes[399], nodes[657],  nodes[1296]);
    tranif1 (nodes[373], nodes[657],  nodes[1453]);
    tranif1 (nodes[264], nodes[558],  nodes[1312]);
    tranif1 (nodes[812], nodes[558],  nodes[646]);
    tranif1 (nodes[210], nodes[1513],  nodes[943]);
    tranif1 (nodes[1706], nodes[1500],  nodes[379]);
    tranif1 (nodes[1345], nodes[558],  nodes[379]);
    tranif1 (nodes[1508], nodes[1101],  nodes[813]);
    tranif1 (nodes[11], nodes[558],  nodes[4]);
    tranif1 (nodes[558], nodes[1380],  nodes[819]);
    tranif1 (nodes[657], nodes[214],  nodes[714]);
    tranif1 (nodes[558], nodes[818],  nodes[43]);
    tranif1 (nodes[1107], nodes[558],  nodes[1520]);
    tranif1 (nodes[1130], nodes[558],  nodes[1002]);
    tranif1 (nodes[805], nodes[779],  nodes[943]);
    tranif1 (nodes[101], nodes[1141],  nodes[710]);
    tranif1 (nodes[1308], nodes[408],  nodes[943]);
    tranif1 (nodes[379], nodes[1480],  nodes[1581]);
    tranif1 (nodes[191], nodes[558],  nodes[347]);
    tranif1 (nodes[558], nodes[1116],  nodes[1537]);
    tranif1 (nodes[1116], nodes[558],  nodes[1537]);
    tranif1 (nodes[558], nodes[1116],  nodes[1537]);
    tranif1 (nodes[558], nodes[169],  nodes[1624]);
    tranif1 (nodes[558], nodes[938],  nodes[408]);
    tranif1 (nodes[558], nodes[1125],  nodes[1576]);
    tranif1 (nodes[1394], nodes[1609],  nodes[943]);
    tranif1 (nodes[558], nodes[453],  nodes[205]);
    tranif1 (nodes[368], nodes[558],  nodes[309]);
    tranif1 (nodes[1172], nodes[405],  nodes[1544]);
    tranif1 (nodes[373], nodes[558],  nodes[1720]);
    tranif1 (nodes[612], nodes[657],  nodes[1720]);
    tranif1 (nodes[657], nodes[1076],  nodes[1088]);
    tranif1 (nodes[773], nodes[558],  nodes[646]);
    tranif1 (nodes[1141], nodes[558],  nodes[982]);
    tranif1 (nodes[1203], nodes[558],  nodes[1135]);
    tranif1 (nodes[1629], nodes[558],  nodes[1135]);
    tranif1 (nodes[813], nodes[558],  nodes[1258]);
    tranif1 (nodes[720], nodes[558],  nodes[248]);
    tranif1 (nodes[1371], nodes[558],  nodes[1045]);
    tranif1 (nodes[1237], nodes[558],  nodes[999]);
    tranif1 (nodes[558], nodes[1237],  nodes[999]);
    tranif1 (nodes[1237], nodes[558],  nodes[999]);
    tranif1 (nodes[1237], nodes[558],  nodes[999]);
    tranif1 (nodes[558], nodes[1237],  nodes[999]);
    tranif1 (nodes[1237], nodes[558],  nodes[999]);
    tranif1 (nodes[558], nodes[1237],  nodes[999]);
    tranif1 (nodes[29], nodes[561],  nodes[943]);
    tranif1 (nodes[876], nodes[558],  nodes[867]);
    tranif1 (nodes[1717], nodes[558],  nodes[1173]);
    tranif1 (nodes[558], nodes[206],  nodes[1146]);
    tranif1 (nodes[1106], nodes[558],  nodes[76]);
    tranif1 (nodes[1033], nodes[558],  nodes[241]);
    tranif1 (nodes[1015], nodes[657],  nodes[241]);
    tranif1 (nodes[886], nodes[975],  nodes[995]);
    tranif1 (nodes[1371], nodes[558],  nodes[201]);
    tranif1 (nodes[272], nodes[558],  nodes[273]);
    tranif1 (nodes[558], nodes[307],  nodes[846]);
    tranif1 (nodes[541], nodes[1183],  nodes[879]);
    tranif1 (nodes[380], nodes[558],  nodes[827]);
    tranif1 (nodes[124], nodes[558],  nodes[1061]);
    tranif1 (nodes[1403], nodes[332],  nodes[654]);
    tranif1 (nodes[657], nodes[1108],  nodes[943]);
    tranif1 (nodes[355], nodes[558],  nodes[621]);
    tranif1 (nodes[251], nodes[558],  nodes[1035]);
    tranif1 (nodes[558], nodes[188],  nodes[1606]);
    tranif1 (nodes[719], nodes[407],  nodes[41]);
    tranif1 (nodes[87], nodes[52],  nodes[41]);
    tranif1 (nodes[1424], nodes[1651],  nodes[41]);
    tranif1 (nodes[1661], nodes[315],  nodes[41]);
    tranif1 (nodes[1095], nodes[1160],  nodes[41]);
    tranif1 (nodes[1387], nodes[483],  nodes[41]);
    tranif1 (nodes[1014], nodes[13],  nodes[41]);
    tranif1 (nodes[1147], nodes[1539],  nodes[41]);
    tranif1 (nodes[689], nodes[558],  nodes[370]);
    tranif1 (nodes[1534], nodes[558],  nodes[805]);
    tranif1 (nodes[1136], nodes[326],  nodes[943]);
    tranif1 (nodes[170], nodes[1117],  nodes[943]);
    tranif1 (nodes[873], nodes[797],  nodes[710]);
    tranif1 (nodes[1087], nodes[558],  nodes[1382]);
    tranif1 (nodes[558], nodes[1178],  nodes[960]);
    tranif1 (nodes[316], nodes[1628],  nodes[977]);
    tranif1 (nodes[143], nodes[558],  nodes[977]);
    tranif1 (nodes[166], nodes[1098],  nodes[874]);
    tranif1 (nodes[1336], nodes[1212],  nodes[874]);
    tranif1 (nodes[1188], nodes[1532],  nodes[874]);
    tranif1 (nodes[1702], nodes[1405],  nodes[874]);
    tranif1 (nodes[1150], nodes[183],  nodes[874]);
    tranif1 (nodes[1287], nodes[81],  nodes[874]);
    tranif1 (nodes[558], nodes[802],  nodes[781]);
    tranif1 (nodes[406], nodes[558],  nodes[1525]);
    tranif1 (nodes[555], nodes[558],  nodes[1525]);
    tranif1 (nodes[558], nodes[427],  nodes[647]);
    tranif1 (nodes[558], nodes[1425],  nodes[1372]);
    tranif1 (nodes[1648], nodes[242],  nodes[943]);
    tranif1 (nodes[1674], nodes[931],  nodes[710]);
    tranif1 (nodes[1450], nodes[1526],  nodes[710]);
    tranif1 (nodes[558], nodes[638],  nodes[1273]);
    tranif1 (nodes[154], nodes[558],  nodes[512]);
    tranif1 (nodes[558], nodes[874],  nodes[1247]);
    tranif1 (nodes[1448], nodes[558],  nodes[1427]);
    tranif1 (nodes[1357], nodes[558],  nodes[223]);
    tranif1 (nodes[1002], nodes[558],  nodes[1219]);
    tranif1 (nodes[687], nodes[1108],  nodes[1042]);
    tranif1 (nodes[1477], nodes[604],  nodes[943]);
    tranif1 (nodes[1082], nodes[367],  nodes[206]);
    tranif1 (nodes[558], nodes[818],  nodes[265]);
    tranif1 (nodes[971], nodes[558],  nodes[1575]);
    tranif1 (nodes[406], nodes[371],  nodes[105]);
    tranif1 (nodes[555], nodes[558],  nodes[105]);
    tranif1 (nodes[1323], nodes[558],  nodes[631]);
    tranif1 (nodes[283], nodes[657],  nodes[631]);
    tranif1 (nodes[558], nodes[267],  nodes[544]);
    tranif1 (nodes[558], nodes[616],  nodes[1482]);
    tranif1 (nodes[1437], nodes[657],  nodes[943]);
    tranif1 (nodes[1364], nodes[558],  nodes[101]);
    tranif1 (nodes[844], nodes[558],  nodes[985]);
    tranif1 (nodes[1151], nodes[558],  nodes[1262]);
    tranif1 (nodes[1212], nodes[618],  nodes[654]);
    tranif1 (nodes[1098], nodes[280],  nodes[654]);
    tranif1 (nodes[1702], nodes[3],  nodes[654]);
    tranif1 (nodes[1532], nodes[998],  nodes[654]);
    tranif1 (nodes[81], nodes[1389],  nodes[654]);
    tranif1 (nodes[183], nodes[694],  nodes[654]);
    tranif1 (nodes[883], nodes[558],  nodes[315]);
    tranif1 (nodes[178], nodes[558],  nodes[1307]);
    tranif1 (nodes[347], nodes[558],  nodes[281]);
    tranif1 (nodes[558], nodes[553],  nodes[781]);
    tranif1 (nodes[1235], nodes[558],  nodes[1413]);
    tranif1 (nodes[1649], nodes[558],  nodes[764]);
    tranif1 (nodes[1187], nodes[558],  nodes[1212]);
    tranif1 (nodes[1597], nodes[719],  nodes[710]);
    tranif1 (nodes[1605], nodes[558],  nodes[1410]);
    tranif1 (nodes[558], nodes[455],  nodes[279]);
    tranif1 (nodes[657], nodes[407],  nodes[943]);
    tranif1 (nodes[558], nodes[1724],  nodes[730]);
    tranif1 (nodes[175], nodes[558],  nodes[612]);
    tranif1 (nodes[175], nodes[558],  nodes[612]);
    tranif1 (nodes[175], nodes[558],  nodes[612]);
    tranif1 (nodes[175], nodes[558],  nodes[612]);
    tranif1 (nodes[558], nodes[175],  nodes[612]);
    tranif1 (nodes[558], nodes[175],  nodes[612]);
    tranif1 (nodes[175], nodes[558],  nodes[612]);
    tranif1 (nodes[317], nodes[558],  nodes[445]);
    tranif1 (nodes[417], nodes[558],  nodes[445]);
    tranif1 (nodes[417], nodes[558],  nodes[445]);
    tranif1 (nodes[558], nodes[127],  nodes[710]);
    tranif1 (nodes[558], nodes[539],  nodes[445]);
    tranif1 (nodes[539], nodes[558],  nodes[445]);
    tranif1 (nodes[558], nodes[539],  nodes[445]);
    tranif1 (nodes[539], nodes[558],  nodes[445]);
    tranif1 (nodes[539], nodes[558],  nodes[445]);
    tranif1 (nodes[558], nodes[287],  nodes[768]);
    tranif1 (nodes[558], nodes[1215],  nodes[1382]);
    tranif1 (nodes[547], nodes[558],  nodes[1220]);
    tranif1 (nodes[558], nodes[817],  nodes[1220]);
    tranif1 (nodes[1242], nodes[1637],  nodes[1015]);
    tranif1 (nodes[872], nodes[1282],  nodes[1015]);
    tranif1 (nodes[401], nodes[413],  nodes[1015]);
    tranif1 (nodes[1464], nodes[558],  nodes[784]);
    tranif1 (nodes[501], nodes[558],  nodes[67]);
    tranif1 (nodes[913], nodes[558],  nodes[1699]);
    tranif1 (nodes[558], nodes[261],  nodes[447]);
    tranif1 (nodes[558], nodes[388],  nodes[425]);
    tranif1 (nodes[54], nodes[564],  nodes[801]);
    tranif1 (nodes[558], nodes[335],  nodes[347]);
    tranif1 (nodes[1596], nodes[558],  nodes[1602]);
    tranif1 (nodes[558], nodes[442],  nodes[182]);
    tranif1 (nodes[798], nodes[657],  nodes[746]);
    tranif1 (nodes[729], nodes[261],  nodes[943]);
    tranif1 (nodes[323], nodes[959],  nodes[710]);
    tranif1 (nodes[1605], nodes[1183],  nodes[710]);
    tranif1 (nodes[793], nodes[1181],  nodes[1595]);
    tranif1 (nodes[558], nodes[488],  nodes[1227]);
    tranif1 (nodes[558], nodes[182],  nodes[0]);
    tranif1 (nodes[558], nodes[861],  nodes[1452]);
    tranif1 (nodes[1000], nodes[558],  nodes[575]);
    tranif1 (nodes[1055], nodes[558],  nodes[1708]);
    tranif1 (nodes[921], nodes[558],  nodes[1305]);
    tranif1 (nodes[558], nodes[800],  nodes[525]);
    tranif1 (nodes[657], nodes[1331],  nodes[525]);
    tranif1 (nodes[558], nodes[80],  nodes[1130]);
    tranif1 (nodes[980], nodes[558],  nodes[1381]);
    tranif1 (nodes[558], nodes[1133],  nodes[328]);
    tranif1 (nodes[194], nodes[558],  nodes[328]);
    tranif1 (nodes[558], nodes[451],  nodes[66]);
    tranif1 (nodes[558], nodes[451],  nodes[66]);
    tranif1 (nodes[558], nodes[451],  nodes[66]);
    tranif1 (nodes[558], nodes[451],  nodes[66]);
    tranif1 (nodes[48], nodes[558],  nodes[943]);
    tranif1 (nodes[741], nodes[558],  nodes[943]);
    tranif1 (nodes[558], nodes[600],  nodes[1341]);
    tranif1 (nodes[300], nodes[558],  nodes[712]);
    tranif1 (nodes[1224], nodes[558],  nodes[1108]);
    tranif1 (nodes[1397], nodes[1303],  nodes[335]);
    tranif1 (nodes[558], nodes[279],  nodes[253]);
    tranif1 (nodes[558], nodes[1692],  nodes[253]);
    tranif1 (nodes[943], nodes[657],  nodes[1129]);
    tranif1 (nodes[558], nodes[906],  nodes[1333]);
    tranif1 (nodes[558], nodes[82],  nodes[558]);
    tranif1 (nodes[605], nodes[558],  nodes[1081]);
    tranif1 (nodes[1198], nodes[558],  nodes[1530]);
    tranif1 (nodes[248], nodes[657],  nodes[424]);
    tranif1 (nodes[1178], nodes[558],  nodes[614]);
    tranif1 (nodes[558], nodes[248],  nodes[198]);
    tranif1 (nodes[558], nodes[424],  nodes[198]);
    tranif1 (nodes[1604], nodes[1717],  nodes[335]);
    tranif1 (nodes[977], nodes[413],  nodes[437]);
    tranif1 (nodes[1054], nodes[558],  nodes[926]);
    tranif1 (nodes[1150], nodes[694],  nodes[1700]);
    tranif1 (nodes[349], nodes[558],  nodes[869]);
    tranif1 (nodes[349], nodes[558],  nodes[869]);
    tranif1 (nodes[558], nodes[349],  nodes[869]);
    tranif1 (nodes[349], nodes[558],  nodes[869]);
    tranif1 (nodes[558], nodes[349],  nodes[869]);
    tranif1 (nodes[558], nodes[349],  nodes[869]);
    tranif1 (nodes[558], nodes[349],  nodes[869]);
    tranif1 (nodes[1393], nodes[657],  nodes[1076]);
    tranif1 (nodes[1393], nodes[657],  nodes[1076]);
    tranif1 (nodes[641], nodes[558],  nodes[1611]);
    tranif1 (nodes[166], nodes[280],  nodes[1700]);
    tranif1 (nodes[544], nodes[558],  nodes[244]);
    tranif1 (nodes[939], nodes[757],  nodes[1144]);
    tranif1 (nodes[428], nodes[1456],  nodes[248]);
    tranif1 (nodes[1091], nodes[12],  nodes[248]);
    tranif1 (nodes[16], nodes[558],  nodes[248]);
    tranif1 (nodes[558], nodes[213],  nodes[82]);
    tranif1 (nodes[686], nodes[558],  nodes[170]);
    tranif1 (nodes[280], nodes[558],  nodes[601]);
    tranif1 (nodes[162], nodes[1654],  nodes[943]);
    tranif1 (nodes[1062], nodes[705],  nodes[821]);
    tranif1 (nodes[558], nodes[6],  nodes[521]);
    tranif1 (nodes[417], nodes[657],  nodes[317]);
    tranif1 (nodes[52], nodes[558],  nodes[203]);
    tranif1 (nodes[1076], nodes[558],  nodes[353]);
    tranif1 (nodes[1076], nodes[558],  nodes[353]);
    tranif1 (nodes[1463], nodes[558],  nodes[353]);
    tranif1 (nodes[845], nodes[1553],  nodes[710]);
    tranif1 (nodes[558], nodes[1358],  nodes[1109]);
    tranif1 (nodes[1281], nodes[558],  nodes[650]);
    tranif1 (nodes[500], nodes[558],  nodes[427]);
    tranif1 (nodes[1314], nodes[112],  nodes[427]);
    tranif1 (nodes[462], nodes[878],  nodes[943]);
    tranif1 (nodes[558], nodes[807],  nodes[330]);
    tranif1 (nodes[1716], nodes[558],  nodes[1258]);
    tranif1 (nodes[315], nodes[584],  nodes[48]);
    tranif1 (nodes[1651], nodes[502],  nodes[48]);
    tranif1 (nodes[483], nodes[49],  nodes[48]);
    tranif1 (nodes[1160], nodes[948],  nodes[48]);
    tranif1 (nodes[1539], nodes[205],  nodes[48]);
    tranif1 (nodes[13], nodes[1551],  nodes[48]);
    tranif1 (nodes[657], nodes[1336],  nodes[943]);
    tranif1 (nodes[1029], nodes[1187],  nodes[943]);
    tranif1 (nodes[1383], nodes[558],  nodes[1503]);
    tranif1 (nodes[92], nodes[1667],  nodes[821]);
    tranif1 (nodes[1683], nodes[1090],  nodes[943]);
    tranif1 (nodes[1018], nodes[558],  nodes[762]);
    tranif1 (nodes[558], nodes[421],  nodes[135]);
    tranif1 (nodes[558], nodes[421],  nodes[135]);
    tranif1 (nodes[421], nodes[558],  nodes[135]);
    tranif1 (nodes[558], nodes[421],  nodes[135]);
    tranif1 (nodes[657], nodes[1160],  nodes[943]);
    tranif1 (nodes[657], nodes[1630],  nodes[943]);
    tranif1 (nodes[1012], nodes[366],  nodes[440]);
    tranif1 (nodes[558], nodes[1143],  nodes[668]);
    tranif1 (nodes[558], nodes[21],  nodes[1162]);
    tranif1 (nodes[15], nodes[474],  nodes[943]);
    tranif1 (nodes[54], nodes[1169],  nodes[1263]);
    tranif1 (nodes[1035], nodes[558],  nodes[962]);
    tranif1 (nodes[558], nodes[963],  nodes[1523]);
    tranif1 (nodes[657], nodes[635],  nodes[1523]);
    tranif1 (nodes[558], nodes[1413],  nodes[1260]);
    tranif1 (nodes[1235], nodes[657],  nodes[1260]);
    tranif1 (nodes[130], nodes[558],  nodes[220]);
    tranif1 (nodes[657], nodes[639],  nodes[220]);
    tranif1 (nodes[102], nodes[558],  nodes[400]);
    tranif1 (nodes[1696], nodes[657],  nodes[400]);
    tranif1 (nodes[1696], nodes[558],  nodes[834]);
    tranif1 (nodes[400], nodes[558],  nodes[834]);
    tranif1 (nodes[558], nodes[1561],  nodes[777]);
    tranif1 (nodes[558], nodes[656],  nodes[604]);
    tranif1 (nodes[657], nodes[1443],  nodes[1545]);
    tranif1 (nodes[1012], nodes[558],  nodes[1246]);
    tranif1 (nodes[949], nodes[558],  nodes[1334]);
    tranif1 (nodes[1406], nodes[558],  nodes[1334]);
    tranif1 (nodes[1108], nodes[977],  nodes[859]);
    tranif1 (nodes[187], nodes[402],  nodes[710]);
    tranif1 (nodes[1129], nodes[558],  nodes[358]);
    tranif1 (nodes[1129], nodes[558],  nodes[358]);
    tranif1 (nodes[1113], nodes[1717],  nodes[943]);
    tranif1 (nodes[1001], nodes[871],  nodes[1263]);
    tranif1 (nodes[52], nodes[657],  nodes[943]);
    tranif1 (nodes[498], nodes[568],  nodes[943]);
    tranif1 (nodes[558], nodes[138],  nodes[1250]);
    tranif1 (nodes[558], nodes[990],  nodes[1250]);
    tranif1 (nodes[657], nodes[1041],  nodes[1250]);
    tranif1 (nodes[1214], nodes[558],  nodes[1011]);
    tranif1 (nodes[182], nodes[558],  nodes[1655]);
    tranif1 (nodes[558], nodes[1356],  nodes[1136]);
    tranif1 (nodes[558], nodes[909],  nodes[378]);
    tranif1 (nodes[558], nodes[71],  nodes[35]);
    tranif1 (nodes[657], nodes[654],  nodes[35]);
    tranif1 (nodes[558], nodes[1180],  nodes[554]);
    tranif1 (nodes[964], nodes[558],  nodes[554]);
    tranif1 (nodes[558], nodes[1304],  nodes[787]);
    tranif1 (nodes[558], nodes[1347],  nodes[967]);
    tranif1 (nodes[104], nodes[558],  nodes[967]);
    tranif1 (nodes[343], nodes[571],  nodes[710]);
    tranif1 (nodes[1061], nodes[207],  nodes[943]);
    tranif1 (nodes[1004], nodes[473],  nodes[980]);
    tranif1 (nodes[958], nodes[558],  nodes[89]);
    tranif1 (nodes[672], nodes[657],  nodes[963]);
    tranif1 (nodes[558], nodes[863],  nodes[1240]);
    tranif1 (nodes[333], nodes[164],  nodes[943]);
    tranif1 (nodes[1197], nodes[558],  nodes[174]);
    tranif1 (nodes[1170], nodes[558],  nodes[781]);
    tranif1 (nodes[657], nodes[1417],  nodes[670]);
    tranif1 (nodes[1443], nodes[558],  nodes[994]);
    tranif1 (nodes[558], nodes[1443],  nodes[994]);
    tranif1 (nodes[1443], nodes[558],  nodes[994]);
    tranif1 (nodes[1443], nodes[558],  nodes[994]);
    tranif1 (nodes[558], nodes[1443],  nodes[994]);
    tranif1 (nodes[1443], nodes[558],  nodes[994]);
    tranif1 (nodes[558], nodes[1443],  nodes[994]);
    tranif1 (nodes[518], nodes[558],  nodes[1439]);
    tranif1 (nodes[721], nodes[1435],  nodes[654]);
    tranif1 (nodes[880], nodes[558],  nodes[13]);
    tranif1 (nodes[558], nodes[747],  nodes[670]);
    tranif1 (nodes[558], nodes[1480],  nodes[1472]);
    tranif1 (nodes[558], nodes[1294],  nodes[1587]);
    tranif1 (nodes[1083], nodes[558],  nodes[1587]);
    tranif1 (nodes[942], nodes[1285],  nodes[1628]);
    tranif1 (nodes[877], nodes[558],  nodes[506]);
    tranif1 (nodes[1642], nodes[1278],  nodes[824]);
    tranif1 (nodes[1084], nodes[722],  nodes[59]);
    tranif1 (nodes[558], nodes[1347],  nodes[1396]);
    tranif1 (nodes[634], nodes[558],  nodes[1676]);
    tranif1 (nodes[657], nodes[86],  nodes[1676]);
    tranif1 (nodes[310], nodes[194],  nodes[943]);
    tranif1 (nodes[558], nodes[1092],  nodes[118]);
    tranif1 (nodes[572], nodes[558],  nodes[1176]);
    tranif1 (nodes[558], nodes[61],  nodes[1336]);
    tranif1 (nodes[558], nodes[268],  nodes[1100]);
    tranif1 (nodes[558], nodes[268],  nodes[1100]);
    tranif1 (nodes[558], nodes[268],  nodes[1100]);
    tranif1 (nodes[383], nodes[558],  nodes[712]);
    tranif1 (nodes[558], nodes[1560],  nodes[1337]);
    tranif1 (nodes[3], nodes[558],  nodes[1603]);
    tranif1 (nodes[754], nodes[1422],  nodes[443]);
    tranif1 (nodes[755], nodes[558],  nodes[443]);
    tranif1 (nodes[601], nodes[496],  nodes[943]);
    tranif1 (nodes[558], nodes[225],  nodes[1223]);
    tranif1 (nodes[859], nodes[657],  nodes[1223]);
    tranif1 (nodes[558], nodes[895],  nodes[337]);
    tranif1 (nodes[1222], nodes[558],  nodes[1225]);
    tranif1 (nodes[870], nodes[87],  nodes[710]);
    tranif1 (nodes[1414], nodes[684],  nodes[1015]);
    tranif1 (nodes[606], nodes[1437],  nodes[1015]);
    tranif1 (nodes[459], nodes[844],  nodes[943]);
    tranif1 (nodes[558], nodes[568],  nodes[175]);
    tranif1 (nodes[558], nodes[916],  nodes[1517]);
    tranif1 (nodes[1299], nodes[765],  nodes[1015]);
    tranif1 (nodes[314], nodes[1630],  nodes[1015]);
    tranif1 (nodes[331], nodes[121],  nodes[1015]);
    tranif1 (nodes[57], nodes[1402],  nodes[293]);
    tranif1 (nodes[356], nodes[207],  nodes[293]);
    tranif1 (nodes[558], nodes[810],  nodes[293]);
    tranif1 (nodes[1106], nodes[734],  nodes[335]);
    tranif1 (nodes[558], nodes[330],  nodes[807]);
    tranif1 (nodes[558], nodes[1041],  nodes[990]);
    tranif1 (nodes[657], nodes[138],  nodes[990]);
    tranif1 (nodes[1575], nodes[558],  nodes[1357]);
    tranif1 (nodes[1475], nodes[558],  nodes[1097]);
    tranif1 (nodes[1691], nodes[740],  nodes[59]);
    tranif1 (nodes[29], nodes[51],  nodes[787]);
    tranif1 (nodes[203], nodes[558],  nodes[1635]);
    tranif1 (nodes[237], nodes[1641],  nodes[710]);
    tranif1 (nodes[409], nodes[724],  nodes[710]);
    tranif1 (nodes[845], nodes[1426],  nodes[1662]);
    tranif1 (nodes[80], nodes[558],  nodes[267]);
    tranif1 (nodes[916], nodes[387],  nodes[206]);
    tranif1 (nodes[1071], nodes[649],  nodes[59]);
    tranif1 (nodes[1572], nodes[22],  nodes[505]);
    tranif1 (nodes[193], nodes[558],  nodes[505]);
    tranif1 (nodes[495], nodes[1071],  nodes[943]);
    tranif1 (nodes[558], nodes[1130],  nodes[1109]);
    tranif1 (nodes[558], nodes[1163],  nodes[1417]);
    tranif1 (nodes[1163], nodes[558],  nodes[1417]);
    tranif1 (nodes[558], nodes[1163],  nodes[1417]);
    tranif1 (nodes[1163], nodes[558],  nodes[1417]);
    tranif1 (nodes[558], nodes[1163],  nodes[1417]);
    tranif1 (nodes[116], nodes[718],  nodes[943]);
    tranif1 (nodes[558], nodes[165],  nodes[1236]);
    tranif1 (nodes[345], nodes[1584],  nodes[8]);
    tranif1 (nodes[37], nodes[558],  nodes[1634]);
    tranif1 (nodes[224], nodes[558],  nodes[1634]);
    tranif1 (nodes[558], nodes[176],  nodes[10]);
    tranif1 (nodes[558], nodes[628],  nodes[55]);
    tranif1 (nodes[1616], nodes[299],  nodes[1614]);
    tranif1 (nodes[335], nodes[558],  nodes[925]);
    tranif1 (nodes[1697], nodes[558],  nodes[664]);
    tranif1 (nodes[1134], nodes[558],  nodes[1465]);
    tranif1 (nodes[558], nodes[122],  nodes[1459]);
    tranif1 (nodes[558], nodes[1030],  nodes[1459]);
    tranif1 (nodes[1305], nodes[558],  nodes[772]);
    tranif1 (nodes[921], nodes[657],  nodes[772]);
    tranif1 (nodes[496], nodes[558],  nodes[1098]);
    tranif1 (nodes[558], nodes[481],  nodes[1079]);
    tranif1 (nodes[558], nodes[534],  nodes[943]);
    tranif1 (nodes[558], nodes[625],  nodes[459]);
    tranif1 (nodes[558], nodes[830],  nodes[43]);
    tranif1 (nodes[558], nodes[103],  nodes[558]);
    tranif1 (nodes[580], nodes[566],  nodes[755]);
    tranif1 (nodes[657], nodes[520],  nodes[1634]);
    tranif1 (nodes[17], nodes[558],  nodes[732]);
    tranif1 (nodes[1536], nodes[558],  nodes[732]);
    tranif1 (nodes[1679], nodes[248],  nodes[710]);
    tranif1 (nodes[1215], nodes[223],  nodes[710]);
    tranif1 (nodes[558], nodes[1327],  nodes[748]);
    tranif1 (nodes[511], nodes[558],  nodes[1078]);
    tranif1 (nodes[719], nodes[1108],  nodes[863]);
    tranif1 (nodes[87], nodes[991],  nodes[863]);
    tranif1 (nodes[1424], nodes[1473],  nodes[863]);
    tranif1 (nodes[1661], nodes[1302],  nodes[863]);
    tranif1 (nodes[1095], nodes[892],  nodes[863]);
    tranif1 (nodes[1387], nodes[1503],  nodes[863]);
    tranif1 (nodes[1014], nodes[833],  nodes[863]);
    tranif1 (nodes[1147], nodes[493],  nodes[863]);
    tranif1 (nodes[558], nodes[1368],  nodes[1374]);
    tranif1 (nodes[1493], nodes[657],  nodes[322]);
    tranif1 (nodes[657], nodes[1493],  nodes[322]);
    tranif1 (nodes[657], nodes[1493],  nodes[322]);
    tranif1 (nodes[657], nodes[1493],  nodes[322]);
    tranif1 (nodes[1233], nodes[558],  nodes[1536]);
    tranif1 (nodes[286], nodes[558],  nodes[1536]);
    tranif1 (nodes[382], nodes[558],  nodes[1536]);
    tranif1 (nodes[1173], nodes[558],  nodes[1536]);
    tranif1 (nodes[1543], nodes[558],  nodes[1536]);
    tranif1 (nodes[76], nodes[558],  nodes[1536]);
    tranif1 (nodes[558], nodes[1658],  nodes[1536]);
    tranif1 (nodes[558], nodes[245],  nodes[1536]);
    tranif1 (nodes[558], nodes[985],  nodes[1536]);
    tranif1 (nodes[682], nodes[558],  nodes[1536]);
    tranif1 (nodes[665], nodes[558],  nodes[1536]);
    tranif1 (nodes[271], nodes[558],  nodes[1536]);
    tranif1 (nodes[552], nodes[558],  nodes[1536]);
    tranif1 (nodes[558], nodes[1623],  nodes[1536]);
    tranif1 (nodes[558], nodes[403],  nodes[1536]);
    tranif1 (nodes[558], nodes[1273],  nodes[1536]);
    tranif1 (nodes[1337], nodes[558],  nodes[1536]);
    tranif1 (nodes[1355], nodes[558],  nodes[1536]);
    tranif1 (nodes[787], nodes[558],  nodes[1536]);
    tranif1 (nodes[575], nodes[558],  nodes[1536]);
    tranif1 (nodes[257], nodes[558],  nodes[1536]);
    tranif1 (nodes[558], nodes[179],  nodes[1536]);
    tranif1 (nodes[558], nodes[131],  nodes[1536]);
    tranif1 (nodes[558], nodes[1420],  nodes[1536]);
    tranif1 (nodes[1342], nodes[558],  nodes[1536]);
    tranif1 (nodes[4], nodes[558],  nodes[1536]);
    tranif1 (nodes[1396], nodes[558],  nodes[1536]);
    tranif1 (nodes[167], nodes[558],  nodes[1536]);
    tranif1 (nodes[303], nodes[558],  nodes[1536]);
    tranif1 (nodes[558], nodes[1504],  nodes[1536]);
    tranif1 (nodes[558], nodes[1721],  nodes[1536]);
    tranif1 (nodes[558], nodes[1074],  nodes[1536]);
    tranif1 (nodes[1478], nodes[558],  nodes[1536]);
    tranif1 (nodes[594], nodes[558],  nodes[1536]);
    tranif1 (nodes[1292], nodes[558],  nodes[1536]);
    tranif1 (nodes[1114], nodes[558],  nodes[1536]);
    tranif1 (nodes[1476], nodes[558],  nodes[1536]);
    tranif1 (nodes[558], nodes[1226],  nodes[1536]);
    tranif1 (nodes[558], nodes[1419],  nodes[1536]);
    tranif1 (nodes[1491], nodes[573],  nodes[943]);
    tranif1 (nodes[272], nodes[558],  nodes[236]);
    tranif1 (nodes[299], nodes[558],  nodes[587]);
    tranif1 (nodes[558], nodes[1466],  nodes[337]);
    tranif1 (nodes[558], nodes[1601],  nodes[337]);
    tranif1 (nodes[1173], nodes[558],  nodes[337]);
    tranif1 (nodes[1562], nodes[558],  nodes[337]);
    tranif1 (nodes[1543], nodes[558],  nodes[337]);
    tranif1 (nodes[1540], nodes[558],  nodes[337]);
    tranif1 (nodes[245], nodes[558],  nodes[337]);
    tranif1 (nodes[558], nodes[985],  nodes[337]);
    tranif1 (nodes[558], nodes[682],  nodes[337]);
    tranif1 (nodes[558], nodes[665],  nodes[337]);
    tranif1 (nodes[286], nodes[558],  nodes[337]);
    tranif1 (nodes[271], nodes[558],  nodes[337]);
    tranif1 (nodes[370], nodes[558],  nodes[337]);
    tranif1 (nodes[403], nodes[558],  nodes[337]);
    tranif1 (nodes[804], nodes[558],  nodes[337]);
    tranif1 (nodes[558], nodes[712],  nodes[337]);
    tranif1 (nodes[558], nodes[546],  nodes[337]);
    tranif1 (nodes[558], nodes[776],  nodes[337]);
    tranif1 (nodes[257], nodes[558],  nodes[337]);
    tranif1 (nodes[179], nodes[558],  nodes[337]);
    tranif1 (nodes[1420], nodes[558],  nodes[337]);
    tranif1 (nodes[4], nodes[558],  nodes[337]);
    tranif1 (nodes[558], nodes[167],  nodes[337]);
    tranif1 (nodes[558], nodes[303],  nodes[337]);
    tranif1 (nodes[558], nodes[1504],  nodes[337]);
    tranif1 (nodes[558], nodes[487],  nodes[337]);
    tranif1 (nodes[579], nodes[558],  nodes[337]);
    tranif1 (nodes[145], nodes[558],  nodes[337]);
    tranif1 (nodes[259], nodes[558],  nodes[337]);
    tranif1 (nodes[517], nodes[558],  nodes[337]);
    tranif1 (nodes[558], nodes[352],  nodes[337]);
    tranif1 (nodes[558], nodes[750],  nodes[337]);
    tranif1 (nodes[558], nodes[528],  nodes[337]);
    tranif1 (nodes[558], nodes[691],  nodes[337]);
    tranif1 (nodes[1646], nodes[558],  nodes[337]);
    tranif1 (nodes[1114], nodes[558],  nodes[337]);
    tranif1 (nodes[1476], nodes[558],  nodes[337]);
    tranif1 (nodes[1226], nodes[558],  nodes[337]);
    tranif1 (nodes[558], nodes[1665],  nodes[337]);
    tranif1 (nodes[558], nodes[840],  nodes[337]);
    tranif1 (nodes[558], nodes[1164],  nodes[337]);
    tranif1 (nodes[848], nodes[473],  nodes[943]);
    tranif1 (nodes[389], nodes[614],  nodes[943]);
    tranif1 (nodes[249], nodes[558],  nodes[1359]);
    tranif1 (nodes[1081], nodes[960],  nodes[943]);
    tranif1 (nodes[558], nodes[1154],  nodes[248]);
    tranif1 (nodes[558], nodes[180],  nodes[248]);
    tranif1 (nodes[1367], nodes[558],  nodes[1202]);
    tranif1 (nodes[57], nodes[558],  nodes[1202]);
    tranif1 (nodes[620], nodes[558],  nodes[307]);
    tranif1 (nodes[256], nodes[558],  nodes[784]);
    tranif1 (nodes[278], nodes[558],  nodes[1551]);
    tranif1 (nodes[558], nodes[171],  nodes[567]);
    tranif1 (nodes[558], nodes[1026],  nodes[567]);
    tranif1 (nodes[322], nodes[657],  nodes[567]);
    tranif1 (nodes[8], nodes[558],  nodes[551]);
    tranif1 (nodes[1125], nodes[1620],  nodes[943]);
    tranif1 (nodes[558], nodes[1297],  nodes[558]);
    tranif1 (nodes[558], nodes[1275],  nodes[832]);
    tranif1 (nodes[558], nodes[437],  nodes[491]);
    tranif1 (nodes[558], nodes[642],  nodes[1502]);
    tranif1 (nodes[558], nodes[951],  nodes[1502]);
    tranif1 (nodes[657], nodes[1152],  nodes[1502]);
    tranif1 (nodes[558], nodes[744],  nodes[892]);
    tranif1 (nodes[696], nodes[911],  nodes[79]);
    tranif1 (nodes[893], nodes[277],  nodes[943]);
    tranif1 (nodes[558], nodes[1257],  nodes[412]);
    tranif1 (nodes[262], nodes[1189],  nodes[1714]);
    tranif1 (nodes[558], nodes[177],  nodes[1241]);
    tranif1 (nodes[351], nodes[558],  nodes[833]);
    tranif1 (nodes[1541], nodes[558],  nodes[43]);
    tranif1 (nodes[91], nodes[558],  nodes[1529]);
    tranif1 (nodes[11], nodes[558],  nodes[167]);
    tranif1 (nodes[1395], nodes[854],  nodes[710]);
    tranif1 (nodes[558], nodes[1290],  nodes[1126]);
    tranif1 (nodes[986], nodes[1556],  nodes[699]);
    tranif1 (nodes[558], nodes[867],  nodes[699]);
    tranif1 (nodes[558], nodes[1649],  nodes[1057]);
    tranif1 (nodes[1538], nodes[558],  nodes[1070]);
    tranif1 (nodes[558], nodes[1334],  nodes[1070]);
    tranif1 (nodes[200], nodes[558],  nodes[1070]);
    tranif1 (nodes[558], nodes[382],  nodes[1112]);
    tranif1 (nodes[558], nodes[1233],  nodes[1112]);
    tranif1 (nodes[558], nodes[84],  nodes[1112]);
    tranif1 (nodes[558], nodes[1543],  nodes[1112]);
    tranif1 (nodes[558], nodes[76],  nodes[1112]);
    tranif1 (nodes[558], nodes[1658],  nodes[1112]);
    tranif1 (nodes[558], nodes[786],  nodes[1112]);
    tranif1 (nodes[558], nodes[1664],  nodes[1112]);
    tranif1 (nodes[558], nodes[1482],  nodes[1112]);
    tranif1 (nodes[558], nodes[286],  nodes[1112]);
    tranif1 (nodes[558], nodes[271],  nodes[1112]);
    tranif1 (nodes[558], nodes[370],  nodes[1112]);
    tranif1 (nodes[558], nodes[552],  nodes[1112]);
    tranif1 (nodes[558], nodes[1612],  nodes[1112]);
    tranif1 (nodes[558], nodes[1487],  nodes[1112]);
    tranif1 (nodes[558], nodes[784],  nodes[1112]);
    tranif1 (nodes[558], nodes[764],  nodes[1112]);
    tranif1 (nodes[558], nodes[1057],  nodes[1112]);
    tranif1 (nodes[558], nodes[1582],  nodes[1112]);
    tranif1 (nodes[558], nodes[1031],  nodes[1112]);
    tranif1 (nodes[558], nodes[804],  nodes[1112]);
    tranif1 (nodes[558], nodes[1311],  nodes[1112]);
    tranif1 (nodes[558], nodes[1428],  nodes[1112]);
    tranif1 (nodes[558], nodes[1520],  nodes[1112]);
    tranif1 (nodes[558], nodes[1259],  nodes[1112]);
    tranif1 (nodes[558], nodes[857],  nodes[1112]);
    tranif1 (nodes[558], nodes[712],  nodes[1112]);
    tranif1 (nodes[558], nodes[1337],  nodes[1112]);
    tranif1 (nodes[558], nodes[1381],  nodes[1112]);
    tranif1 (nodes[558], nodes[776],  nodes[1112]);
    tranif1 (nodes[558], nodes[157],  nodes[1112]);
    tranif1 (nodes[558], nodes[1324],  nodes[1112]);
    tranif1 (nodes[558], nodes[179],  nodes[1112]);
    tranif1 (nodes[558], nodes[131],  nodes[1112]);
    tranif1 (nodes[558], nodes[4],  nodes[1112]);
    tranif1 (nodes[558], nodes[1396],  nodes[1112]);
    tranif1 (nodes[558], nodes[167],  nodes[1112]);
    tranif1 (nodes[558], nodes[303],  nodes[1112]);
    tranif1 (nodes[558], nodes[1086],  nodes[1112]);
    tranif1 (nodes[558], nodes[1074],  nodes[1112]);
    tranif1 (nodes[558], nodes[487],  nodes[1112]);
    tranif1 (nodes[558], nodes[579],  nodes[1112]);
    tranif1 (nodes[558], nodes[0],  nodes[1112]);
    tranif1 (nodes[558], nodes[1478],  nodes[1112]);
    tranif1 (nodes[558], nodes[594],  nodes[1112]);
    tranif1 (nodes[558], nodes[1210],  nodes[1112]);
    tranif1 (nodes[558], nodes[1557],  nodes[1112]);
    tranif1 (nodes[558], nodes[259],  nodes[1112]);
    tranif1 (nodes[558], nodes[1052],  nodes[1112]);
    tranif1 (nodes[558], nodes[791],  nodes[1112]);
    tranif1 (nodes[558], nodes[352],  nodes[1112]);
    tranif1 (nodes[558], nodes[750],  nodes[1112]);
    tranif1 (nodes[558], nodes[932],  nodes[1112]);
    tranif1 (nodes[558], nodes[1589],  nodes[1112]);
    tranif1 (nodes[558], nodes[446],  nodes[1112]);
    tranif1 (nodes[558], nodes[528],  nodes[1112]);
    tranif1 (nodes[558], nodes[309],  nodes[1112]);
    tranif1 (nodes[558], nodes[1430],  nodes[1112]);
    tranif1 (nodes[558], nodes[1646],  nodes[1112]);
    tranif1 (nodes[558], nodes[1476],  nodes[1112]);
    tranif1 (nodes[558], nodes[1226],  nodes[1112]);
    tranif1 (nodes[558], nodes[1569],  nodes[1112]);
    tranif1 (nodes[558], nodes[950],  nodes[1112]);
    tranif1 (nodes[558], nodes[1665],  nodes[1112]);
    tranif1 (nodes[558], nodes[1710],  nodes[1112]);
    tranif1 (nodes[558], nodes[1050],  nodes[1112]);
    tranif1 (nodes[558], nodes[607],  nodes[1112]);
    tranif1 (nodes[558], nodes[219],  nodes[1112]);
    tranif1 (nodes[558], nodes[1384],  nodes[1300]);
    tranif1 (nodes[1016], nodes[416],  nodes[710]);
    tranif1 (nodes[1637], nodes[558],  nodes[276]);
    tranif1 (nodes[1330], nodes[586],  nodes[1544]);
    tranif1 (nodes[1330], nodes[586],  nodes[1544]);
    tranif1 (nodes[318], nodes[1607],  nodes[943]);
    tranif1 (nodes[1466], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[271],  nodes[1328]);
    tranif1 (nodes[558], nodes[370],  nodes[1328]);
    tranif1 (nodes[552], nodes[558],  nodes[1328]);
    tranif1 (nodes[1612], nodes[558],  nodes[1328]);
    tranif1 (nodes[1487], nodes[558],  nodes[1328]);
    tranif1 (nodes[784], nodes[558],  nodes[1328]);
    tranif1 (nodes[244], nodes[558],  nodes[1328]);
    tranif1 (nodes[1623], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[764],  nodes[1328]);
    tranif1 (nodes[558], nodes[403],  nodes[1328]);
    tranif1 (nodes[1582], nodes[558],  nodes[1328]);
    tranif1 (nodes[1031], nodes[558],  nodes[1328]);
    tranif1 (nodes[804], nodes[558],  nodes[1328]);
    tranif1 (nodes[1311], nodes[558],  nodes[1328]);
    tranif1 (nodes[1520], nodes[558],  nodes[1328]);
    tranif1 (nodes[857], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[712],  nodes[1328]);
    tranif1 (nodes[1381], nodes[558],  nodes[1328]);
    tranif1 (nodes[546], nodes[558],  nodes[1328]);
    tranif1 (nodes[776], nodes[558],  nodes[1328]);
    tranif1 (nodes[157], nodes[558],  nodes[1328]);
    tranif1 (nodes[1243], nodes[558],  nodes[1328]);
    tranif1 (nodes[1324], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[131],  nodes[1328]);
    tranif1 (nodes[558], nodes[1396],  nodes[1328]);
    tranif1 (nodes[303], nodes[558],  nodes[1328]);
    tranif1 (nodes[1504], nodes[558],  nodes[1328]);
    tranif1 (nodes[1086], nodes[558],  nodes[1328]);
    tranif1 (nodes[1074], nodes[558],  nodes[1328]);
    tranif1 (nodes[1246], nodes[558],  nodes[1328]);
    tranif1 (nodes[487], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[579],  nodes[1328]);
    tranif1 (nodes[558], nodes[0],  nodes[1328]);
    tranif1 (nodes[1478], nodes[558],  nodes[1328]);
    tranif1 (nodes[594], nodes[558],  nodes[1328]);
    tranif1 (nodes[1557], nodes[558],  nodes[1328]);
    tranif1 (nodes[259], nodes[558],  nodes[1328]);
    tranif1 (nodes[1052], nodes[558],  nodes[1328]);
    tranif1 (nodes[791], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[352],  nodes[1328]);
    tranif1 (nodes[558], nodes[750],  nodes[1328]);
    tranif1 (nodes[932], nodes[558],  nodes[1328]);
    tranif1 (nodes[1589], nodes[558],  nodes[1328]);
    tranif1 (nodes[446], nodes[558],  nodes[1328]);
    tranif1 (nodes[528], nodes[558],  nodes[1328]);
    tranif1 (nodes[309], nodes[558],  nodes[1328]);
    tranif1 (nodes[1430], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[691],  nodes[1328]);
    tranif1 (nodes[558], nodes[1292],  nodes[1328]);
    tranif1 (nodes[1646], nodes[558],  nodes[1328]);
    tranif1 (nodes[1114], nodes[558],  nodes[1328]);
    tranif1 (nodes[1476], nodes[558],  nodes[1328]);
    tranif1 (nodes[1226], nodes[558],  nodes[1328]);
    tranif1 (nodes[1569], nodes[558],  nodes[1328]);
    tranif1 (nodes[1665], nodes[558],  nodes[1328]);
    tranif1 (nodes[558], nodes[1050],  nodes[1328]);
    tranif1 (nodes[1174], nodes[558],  nodes[1328]);
    tranif1 (nodes[1310], nodes[558],  nodes[1063]);
    tranif1 (nodes[657], nodes[672],  nodes[963]);
    tranif1 (nodes[846], nodes[558],  nodes[840]);
    tranif1 (nodes[187], nodes[558],  nodes[1131]);
    tranif1 (nodes[802], nodes[566],  nodes[243]);
    tranif1 (nodes[558], nodes[516],  nodes[216]);
    tranif1 (nodes[558], nodes[1610],  nodes[216]);
    tranif1 (nodes[1046], nodes[558],  nodes[1299]);
    tranif1 (nodes[558], nodes[389],  nodes[1107]);
    tranif1 (nodes[107], nodes[416],  nodes[639]);
    tranif1 (nodes[1334], nodes[558],  nodes[1007]);
    tranif1 (nodes[754], nodes[558],  nodes[1673]);
    tranif1 (nodes[707], nodes[1636],  nodes[639]);
    tranif1 (nodes[558], nodes[1484],  nodes[573]);
    tranif1 (nodes[1013], nodes[558],  nodes[1241]);
    tranif1 (nodes[1217], nodes[558],  nodes[1241]);
    tranif1 (nodes[1157], nodes[558],  nodes[291]);
    tranif1 (nodes[1564], nodes[657],  nodes[291]);
    tranif1 (nodes[558], nodes[1225],  nodes[1524]);
    tranif1 (nodes[10], nodes[558],  nodes[1721]);
    tranif1 (nodes[1488], nodes[558],  nodes[278]);
    tranif1 (nodes[1278], nodes[558],  nodes[462]);
    tranif1 (nodes[558], nodes[725],  nodes[599]);
    tranif1 (nodes[558], nodes[441],  nodes[692]);
    tranif1 (nodes[657], nodes[325],  nodes[692]);
    tranif1 (nodes[300], nodes[558],  nodes[1259]);
    tranif1 (nodes[558], nodes[1350],  nodes[760]);
    tranif1 (nodes[458], nodes[558],  nodes[1473]);
    tranif1 (nodes[558], nodes[27],  nodes[820]);
    tranif1 (nodes[558], nodes[917],  nodes[383]);
    tranif1 (nodes[386], nodes[558],  nodes[622]);
    tranif1 (nodes[558], nodes[1649],  nodes[248]);
    tranif1 (nodes[1366], nodes[472],  nodes[16]);
    tranif1 (nodes[850], nodes[558],  nodes[899]);
    tranif1 (nodes[147], nodes[558],  nodes[353]);
    tranif1 (nodes[147], nodes[558],  nodes[353]);
    tranif1 (nodes[347], nodes[558],  nodes[1385]);
    tranif1 (nodes[1087], nodes[1132],  nodes[710]);
    tranif1 (nodes[558], nodes[1180],  nodes[248]);
    tranif1 (nodes[188], nodes[1373],  nodes[943]);
    tranif1 (nodes[558], nodes[486],  nodes[817]);
    tranif1 (nodes[963], nodes[657],  nodes[997]);
    tranif1 (nodes[558], nodes[1523],  nodes[997]);
    tranif1 (nodes[558], nodes[635],  nodes[997]);
    tranif1 (nodes[558], nodes[859],  nodes[225]);
    tranif1 (nodes[558], nodes[136],  nodes[640]);
    tranif1 (nodes[558], nodes[860],  nodes[640]);
    tranif1 (nodes[558], nodes[1021],  nodes[155]);
    tranif1 (nodes[558], nodes[425],  nodes[155]);
    tranif1 (nodes[1555], nodes[558],  nodes[440]);
    tranif1 (nodes[558], nodes[1686],  nodes[432]);
    tranif1 (nodes[558], nodes[1097],  nodes[432]);
    tranif1 (nodes[672], nodes[558],  nodes[635]);
    tranif1 (nodes[558], nodes[672],  nodes[635]);
    tranif1 (nodes[672], nodes[558],  nodes[635]);
    tranif1 (nodes[558], nodes[672],  nodes[635]);
    tranif1 (nodes[672], nodes[558],  nodes[635]);
    tranif1 (nodes[558], nodes[672],  nodes[635]);
    tranif1 (nodes[558], nodes[672],  nodes[635]);
    tranif1 (nodes[1534], nodes[558],  nodes[43]);
    tranif1 (nodes[558], nodes[1330],  nodes[967]);
    tranif1 (nodes[558], nodes[721],  nodes[181]);
    tranif1 (nodes[683], nodes[1225],  nodes[943]);
    tranif1 (nodes[630], nodes[558],  nodes[726]);
    tranif1 (nodes[1191], nodes[558],  nodes[1195]);
    tranif1 (nodes[657], nodes[1254],  nodes[1195]);
    tranif1 (nodes[558], nodes[1055],  nodes[771]);
    tranif1 (nodes[558], nodes[251],  nodes[221]);
    tranif1 (nodes[251], nodes[558],  nodes[221]);
    tranif1 (nodes[372], nodes[558],  nodes[248]);
    tranif1 (nodes[1085], nodes[1365],  nodes[248]);
    tranif1 (nodes[92], nodes[359],  nodes[943]);
    tranif1 (nodes[756], nodes[626],  nodes[710]);
    tranif1 (nodes[823], nodes[457],  nodes[710]);
    tranif1 (nodes[741], nodes[558],  nodes[255]);
    tranif1 (nodes[657], nodes[148],  nodes[1140]);
    tranif1 (nodes[558], nodes[1634],  nodes[1288]);
    tranif1 (nodes[1040], nodes[558],  nodes[383]);
    tranif1 (nodes[558], nodes[1040],  nodes[383]);
    tranif1 (nodes[699], nodes[558],  nodes[1637]);
    tranif1 (nodes[1495], nodes[1445],  nodes[270]);
    tranif1 (nodes[1552], nodes[558],  nodes[1593]);
    tranif1 (nodes[657], nodes[362],  nodes[1593]);
    tranif1 (nodes[957], nodes[1525],  nodes[1666]);
    tranif1 (nodes[953], nodes[250],  nodes[1666]);
    tranif1 (nodes[740], nodes[701],  nodes[1666]);
    tranif1 (nodes[1071], nodes[884],  nodes[1666]);
    tranif1 (nodes[296], nodes[308],  nodes[1666]);
    tranif1 (nodes[277], nodes[1469],  nodes[1666]);
    tranif1 (nodes[722], nodes[1459],  nodes[1666]);
    tranif1 (nodes[177], nodes[304],  nodes[1666]);
    tranif1 (nodes[256], nodes[558],  nodes[341]);
    tranif1 (nodes[428], nodes[1558],  nodes[16]);
    tranif1 (nodes[591], nodes[252],  nodes[691]);
    tranif1 (nodes[1672], nodes[558],  nodes[558]);
    tranif1 (nodes[558], nodes[1053],  nodes[439]);
    tranif1 (nodes[786], nodes[558],  nodes[156]);
    tranif1 (nodes[1664], nodes[558],  nodes[156]);
    tranif1 (nodes[1482], nodes[558],  nodes[156]);
    tranif1 (nodes[1243], nodes[558],  nodes[156]);
    tranif1 (nodes[822], nodes[558],  nodes[156]);
    tranif1 (nodes[558], nodes[1324],  nodes[156]);
    tranif1 (nodes[1646], nodes[558],  nodes[156]);
    tranif1 (nodes[558], nodes[1155],  nodes[156]);
    tranif1 (nodes[301], nodes[558],  nodes[156]);
    tranif1 (nodes[950], nodes[558],  nodes[156]);
    tranif1 (nodes[1665], nodes[558],  nodes[156]);
    tranif1 (nodes[1710], nodes[558],  nodes[156]);
    tranif1 (nodes[657], nodes[1302],  nodes[943]);
    tranif1 (nodes[1], nodes[1694],  nodes[943]);
    tranif1 (nodes[1403], nodes[54],  nodes[874]);
    tranif1 (nodes[137], nodes[558],  nodes[1120]);
    tranif1 (nodes[558], nodes[1171],  nodes[558]);
    tranif1 (nodes[558], nodes[744],  nodes[833]);
    tranif1 (nodes[558], nodes[218],  nodes[368]);
    tranif1 (nodes[1707], nodes[319],  nodes[623]);
    tranif1 (nodes[558], nodes[388],  nodes[623]);
    tranif1 (nodes[558], nodes[1368],  nodes[1578]);
    tranif1 (nodes[476], nodes[558],  nodes[1027]);
    tranif1 (nodes[558], nodes[368],  nodes[1589]);
    tranif1 (nodes[558], nodes[104],  nodes[1589]);
    tranif1 (nodes[1096], nodes[558],  nodes[153]);
    tranif1 (nodes[558], nodes[1352],  nodes[440]);
    tranif1 (nodes[558], nodes[104],  nodes[440]);
    tranif1 (nodes[558], nodes[812],  nodes[440]);
    tranif1 (nodes[962], nodes[558],  nodes[1585]);
    tranif1 (nodes[558], nodes[1489],  nodes[1398]);
    tranif1 (nodes[1106], nodes[1103],  nodes[258]);
    tranif1 (nodes[558], nodes[1347],  nodes[979]);
    tranif1 (nodes[1464], nodes[558],  nodes[370]);
    tranif1 (nodes[1671], nodes[558],  nodes[955]);
    tranif1 (nodes[558], nodes[911],  nodes[1343]);
    tranif1 (nodes[434], nodes[558],  nodes[790]);
    tranif1 (nodes[70], nodes[558],  nodes[1054]);
    tranif1 (nodes[1106], nodes[558],  nodes[1543]);
    tranif1 (nodes[558], nodes[320],  nodes[1150]);
    tranif1 (nodes[488], nodes[1108],  nodes[283]);
    tranif1 (nodes[1608], nodes[657],  nodes[775]);
    tranif1 (nodes[558], nodes[1423],  nodes[775]);
    tranif1 (nodes[558], nodes[869],  nodes[775]);
    tranif1 (nodes[481], nodes[1473],  nodes[283]);
    tranif1 (nodes[558], nodes[340],  nodes[1164]);
    tranif1 (nodes[1382], nodes[558],  nodes[248]);
    tranif1 (nodes[1053], nodes[673],  nodes[575]);
    tranif1 (nodes[927], nodes[703],  nodes[879]);
    tranif1 (nodes[558], nodes[931],  nodes[415]);
    tranif1 (nodes[558], nodes[1375],  nodes[88]);
    tranif1 (nodes[558], nodes[771],  nodes[1110]);
    tranif1 (nodes[1388], nodes[965],  nodes[1506]);
    tranif1 (nodes[558], nodes[295],  nodes[1506]);
    tranif1 (nodes[7], nodes[558],  nodes[353]);
    tranif1 (nodes[7], nodes[558],  nodes[353]);
    tranif1 (nodes[466], nodes[558],  nodes[353]);
    tranif1 (nodes[558], nodes[920],  nodes[73]);
    tranif1 (nodes[558], nodes[651],  nodes[65]);
    tranif1 (nodes[902], nodes[248],  nodes[710]);
    tranif1 (nodes[558], nodes[1182],  nodes[1384]);
    tranif1 (nodes[895], nodes[1675],  nodes[943]);
    tranif1 (nodes[558], nodes[674],  nodes[25]);
    tranif1 (nodes[829], nodes[1588],  nodes[943]);
    tranif1 (nodes[1281], nodes[894],  nodes[943]);
    tranif1 (nodes[1075], nodes[369],  nodes[943]);
    tranif1 (nodes[1234], nodes[929],  nodes[943]);
    tranif1 (nodes[1223], nodes[558],  nodes[688]);
    tranif1 (nodes[1537], nodes[1638],  nodes[943]);
    tranif1 (nodes[716], nodes[701],  nodes[110]);
    tranif1 (nodes[558], nodes[1716],  nodes[510]);
    tranif1 (nodes[558], nodes[161],  nodes[1113]);
    tranif1 (nodes[558], nodes[1382],  nodes[861]);
    tranif1 (nodes[1068], nodes[558],  nodes[1247]);
    tranif1 (nodes[1591], nodes[1591],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[1591], nodes[558],  nodes[471]);
    tranif1 (nodes[558], nodes[1591],  nodes[471]);
    tranif1 (nodes[1325], nodes[558],  nodes[353]);
    tranif1 (nodes[1325], nodes[558],  nodes[353]);
    tranif1 (nodes[769], nodes[558],  nodes[353]);
    tranif1 (nodes[657], nodes[1467],  nodes[358]);
    tranif1 (nodes[1094], nodes[463],  nodes[710]);
    tranif1 (nodes[1620], nodes[1590],  nodes[879]);
    tranif1 (nodes[1368], nodes[558],  nodes[645]);
    tranif1 (nodes[1275], nodes[558],  nodes[248]);
    tranif1 (nodes[1267], nodes[558],  nodes[52]);
    tranif1 (nodes[514], nodes[494],  nodes[710]);
    tranif1 (nodes[558], nodes[279],  nodes[954]);
    tranif1 (nodes[558], nodes[367],  nodes[954]);
    tranif1 (nodes[1427], nodes[558],  nodes[236]);
    tranif1 (nodes[1464], nodes[558],  nodes[271]);
    tranif1 (nodes[1496], nodes[558],  nodes[114]);
    tranif1 (nodes[843], nodes[1251],  nodes[943]);
    tranif1 (nodes[1519], nodes[558],  nodes[1437]);
    tranif1 (nodes[1447], nodes[262],  nodes[710]);
    tranif1 (nodes[1196], nodes[558],  nodes[522]);
    tranif1 (nodes[153], nodes[246],  nodes[639]);
    tranif1 (nodes[790], nodes[558],  nodes[691]);
    tranif1 (nodes[558], nodes[1601],  nodes[1182]);
    tranif1 (nodes[558], nodes[258],  nodes[1182]);
    tranif1 (nodes[558], nodes[665],  nodes[1182]);
    tranif1 (nodes[558], nodes[764],  nodes[1182]);
    tranif1 (nodes[558], nodes[1057],  nodes[1182]);
    tranif1 (nodes[558], nodes[1381],  nodes[1182]);
    tranif1 (nodes[558], nodes[303],  nodes[1182]);
    tranif1 (nodes[558], nodes[285],  nodes[1182]);
    tranif1 (nodes[558], nodes[594],  nodes[1182]);
    tranif1 (nodes[558], nodes[1052],  nodes[1182]);
    tranif1 (nodes[558], nodes[1589],  nodes[1182]);
    tranif1 (nodes[558], nodes[309],  nodes[1182]);
    tranif1 (nodes[558], nodes[1646],  nodes[1182]);
    tranif1 (nodes[558], nodes[904],  nodes[1182]);
    tranif1 (nodes[558], nodes[1476],  nodes[1182]);
    tranif1 (nodes[558], nodes[950],  nodes[1182]);
    tranif1 (nodes[607], nodes[558],  nodes[1182]);
    tranif1 (nodes[558], nodes[219],  nodes[1182]);
    tranif1 (nodes[984], nodes[558],  nodes[943]);
    tranif1 (nodes[549], nodes[558],  nodes[943]);
    tranif1 (nodes[437], nodes[558],  nodes[943]);
    tranif1 (nodes[859], nodes[558],  nodes[943]);
    tranif1 (nodes[1068], nodes[558],  nodes[943]);
    tranif1 (nodes[654], nodes[558],  nodes[943]);
    tranif1 (nodes[558], nodes[874],  nodes[943]);
    tranif1 (nodes[1167], nodes[558],  nodes[984]);
    tranif1 (nodes[792], nodes[851],  nodes[710]);
    tranif1 (nodes[1248], nodes[558],  nodes[984]);
    tranif1 (nodes[1142], nodes[558],  nodes[984]);
    tranif1 (nodes[1627], nodes[558],  nodes[984]);
    tranif1 (nodes[530], nodes[558],  nodes[984]);
    tranif1 (nodes[510], nodes[558],  nodes[1052]);
    tranif1 (nodes[134], nodes[558],  nodes[1052]);
    tranif1 (nodes[558], nodes[105],  nodes[1165]);
    tranif1 (nodes[942], nodes[558],  nodes[1165]);
    tranif1 (nodes[945], nodes[945],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[945], nodes[558],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[558], nodes[945],  nodes[37]);
    tranif1 (nodes[945], nodes[558],  nodes[37]);
    tranif1 (nodes[558], nodes[36],  nodes[8]);
    tranif1 (nodes[558], nodes[150],  nodes[8]);
    tranif1 (nodes[333], nodes[1030],  nodes[570]);
    tranif1 (nodes[558], nodes[591],  nodes[1258]);
    tranif1 (nodes[657], nodes[684],  nodes[943]);
    tranif1 (nodes[1649], nodes[558],  nodes[1259]);
    tranif1 (nodes[448], nodes[1724],  nodes[943]);
    tranif1 (nodes[1598], nodes[558],  nodes[685]);
    tranif1 (nodes[1060], nodes[558],  nodes[1238]);
    tranif1 (nodes[957], nodes[371],  nodes[921]);
    tranif1 (nodes[250], nodes[965],  nodes[921]);
    tranif1 (nodes[740], nodes[22],  nodes[921]);
    tranif1 (nodes[1071], nodes[274],  nodes[921]);
    tranif1 (nodes[296], nodes[651],  nodes[921]);
    tranif1 (nodes[277], nodes[486],  nodes[921]);
    tranif1 (nodes[1197], nodes[722],  nodes[921]);
    tranif1 (nodes[532], nodes[304],  nodes[921]);
    tranif1 (nodes[1288], nodes[1376],  nodes[710]);
    tranif1 (nodes[327], nodes[558],  nodes[1569]);
    tranif1 (nodes[558], nodes[640],  nodes[988]);
    tranif1 (nodes[828], nodes[34],  nodes[943]);
    tranif1 (nodes[1188], nodes[657],  nodes[943]);
    tranif1 (nodes[2], nodes[558],  nodes[151]);
    tranif1 (nodes[558], nodes[72],  nodes[1326]);
    tranif1 (nodes[597], nodes[1339],  nodes[710]);
    tranif1 (nodes[834], nodes[558],  nodes[402]);
    tranif1 (nodes[558], nodes[436],  nodes[485]);
    tranif1 (nodes[558], nodes[809],  nodes[361]);
    tranif1 (nodes[509], nodes[442],  nodes[943]);
    tranif1 (nodes[564], nodes[558],  nodes[1025]);
    tranif1 (nodes[1601], nodes[558],  nodes[1320]);
    tranif1 (nodes[382], nodes[558],  nodes[1320]);
    tranif1 (nodes[1173], nodes[558],  nodes[1320]);
    tranif1 (nodes[1233], nodes[558],  nodes[1320]);
    tranif1 (nodes[558], nodes[1562],  nodes[1320]);
    tranif1 (nodes[1543], nodes[558],  nodes[1320]);
    tranif1 (nodes[76], nodes[558],  nodes[1320]);
    tranif1 (nodes[1658], nodes[558],  nodes[1320]);
    tranif1 (nodes[1540], nodes[558],  nodes[1320]);
    tranif1 (nodes[245], nodes[558],  nodes[1320]);
    tranif1 (nodes[985], nodes[558],  nodes[1320]);
    tranif1 (nodes[786], nodes[558],  nodes[1320]);
    tranif1 (nodes[558], nodes[1664],  nodes[1320]);
    tranif1 (nodes[682], nodes[558],  nodes[1320]);
    tranif1 (nodes[1482], nodes[558],  nodes[1320]);
    tranif1 (nodes[665], nodes[558],  nodes[1320]);
    tranif1 (nodes[286], nodes[558],  nodes[1320]);
    tranif1 (nodes[324], nodes[558],  nodes[1320]);
    tranif1 (nodes[1337], nodes[558],  nodes[1320]);
    tranif1 (nodes[1355], nodes[558],  nodes[1320]);
    tranif1 (nodes[787], nodes[558],  nodes[1320]);
    tranif1 (nodes[257], nodes[558],  nodes[1320]);
    tranif1 (nodes[179], nodes[558],  nodes[1320]);
    tranif1 (nodes[1420], nodes[558],  nodes[1320]);
    tranif1 (nodes[4], nodes[558],  nodes[1320]);
    tranif1 (nodes[167], nodes[558],  nodes[1320]);
    tranif1 (nodes[145], nodes[558],  nodes[1320]);
    tranif1 (nodes[517], nodes[558],  nodes[1320]);
    tranif1 (nodes[301], nodes[558],  nodes[1320]);
    tranif1 (nodes[950], nodes[558],  nodes[1320]);
    tranif1 (nodes[558], nodes[1710],  nodes[1320]);
    tranif1 (nodes[558], nodes[1419],  nodes[1320]);
    tranif1 (nodes[1164], nodes[558],  nodes[1320]);
    tranif1 (nodes[624], nodes[977],  nodes[1068]);
    tranif1 (nodes[79], nodes[558],  nodes[236]);
    tranif1 (nodes[558], nodes[1003],  nodes[1023]);
    tranif1 (nodes[924], nodes[1425],  nodes[1023]);
    tranif1 (nodes[478], nodes[1645],  nodes[1068]);
    tranif1 (nodes[458], nodes[704],  nodes[1068]);
    tranif1 (nodes[558], nodes[753],  nodes[811]);
    tranif1 (nodes[558], nodes[753],  nodes[811]);
    tranif1 (nodes[127], nodes[558],  nodes[519]);
    tranif1 (nodes[657], nodes[135],  nodes[519]);
    tranif1 (nodes[558], nodes[1575],  nodes[1360]);
    tranif1 (nodes[252], nodes[558],  nodes[1155]);
    tranif1 (nodes[558], nodes[1348],  nodes[1628]);
    tranif1 (nodes[468], nodes[1703],  nodes[16]);
    tranif1 (nodes[558], nodes[366],  nodes[1074]);
    tranif1 (nodes[1583], nodes[308],  nodes[1063]);
    tranif1 (nodes[234], nodes[558],  nodes[1513]);
    tranif1 (nodes[384], nodes[558],  nodes[946]);
    tranif1 (nodes[128], nodes[558],  nodes[1653]);
    tranif1 (nodes[558], nodes[275],  nodes[773]);
    tranif1 (nodes[558], nodes[66],  nodes[376]);
    tranif1 (nodes[842], nodes[558],  nodes[376]);
    tranif1 (nodes[657], nodes[1479],  nodes[376]);
    tranif1 (nodes[1709], nodes[98],  nodes[943]);
    tranif1 (nodes[1282], nodes[558],  nodes[686]);
    tranif1 (nodes[645], nodes[562],  nodes[710]);
    tranif1 (nodes[558], nodes[1705],  nodes[467]);
    tranif1 (nodes[346], nodes[297],  nodes[1392]);
    tranif1 (nodes[284], nodes[558],  nodes[1392]);
    tranif1 (nodes[1227], nodes[558],  nodes[526]);
    tranif1 (nodes[1464], nodes[558],  nodes[552]);
    tranif1 (nodes[78], nodes[558],  nodes[1425]);
    tranif1 (nodes[142], nodes[1310],  nodes[1425]);
    tranif1 (nodes[1617], nodes[558],  nodes[117]);
    tranif1 (nodes[558], nodes[422],  nodes[92]);
    tranif1 (nodes[744], nodes[558],  nodes[991]);
    tranif1 (nodes[558], nodes[851],  nodes[1294]);
    tranif1 (nodes[944], nodes[197],  nodes[943]);
    tranif1 (nodes[1106], nodes[558],  nodes[1658]);
    tranif1 (nodes[1418], nodes[1684],  nodes[710]);
    tranif1 (nodes[558], nodes[388],  nodes[516]);
    tranif1 (nodes[558], nodes[1566],  nodes[1221]);
    tranif1 (nodes[1044], nodes[558],  nodes[812]);
    tranif1 (nodes[1131], nodes[1352],  nodes[943]);
    tranif1 (nodes[1560], nodes[558],  nodes[1355]);
    tranif1 (nodes[95], nodes[1375],  nodes[710]);
    tranif1 (nodes[1529], nodes[1089],  nodes[710]);
    tranif1 (nodes[946], nodes[454],  nodes[844]);
    tranif1 (nodes[1336], nodes[331],  nodes[129]);
    tranif1 (nodes[166], nodes[314],  nodes[129]);
    tranif1 (nodes[606], nodes[1405],  nodes[129]);
    tranif1 (nodes[1188], nodes[1414],  nodes[129]);
    tranif1 (nodes[558], nodes[1391],  nodes[352]);
    tranif1 (nodes[558], nodes[1352],  nodes[352]);
    tranif1 (nodes[1657], nodes[820],  nodes[943]);
    tranif1 (nodes[845], nodes[511],  nodes[553]);
    tranif1 (nodes[608], nodes[558],  nodes[1272]);
    tranif1 (nodes[123], nodes[558],  nodes[413]);
    tranif1 (nodes[185], nodes[558],  nodes[1142]);
    tranif1 (nodes[404], nodes[558],  nodes[1142]);
    tranif1 (nodes[558], nodes[21],  nodes[43]);
    tranif1 (nodes[944], nodes[558],  nodes[1449]);
    tranif1 (nodes[558], nodes[337],  nodes[1675]);
    tranif1 (nodes[1091], nodes[363],  nodes[16]);
    tranif1 (nodes[1717], nodes[558],  nodes[1233]);
    tranif1 (nodes[558], nodes[885],  nodes[384]);
    tranif1 (nodes[558], nodes[550],  nodes[384]);
    tranif1 (nodes[598], nodes[176],  nodes[943]);
    tranif1 (nodes[1653], nodes[1592],  nodes[943]);
    tranif1 (nodes[891], nodes[558],  nodes[943]);
    tranif1 (nodes[1562], nodes[558],  nodes[702]);
    tranif1 (nodes[558], nodes[1543],  nodes[702]);
    tranif1 (nodes[558], nodes[76],  nodes[702]);
    tranif1 (nodes[558], nodes[1540],  nodes[702]);
    tranif1 (nodes[558], nodes[245],  nodes[702]);
    tranif1 (nodes[558], nodes[985],  nodes[702]);
    tranif1 (nodes[558], nodes[786],  nodes[702]);
    tranif1 (nodes[558], nodes[682],  nodes[702]);
    tranif1 (nodes[558], nodes[244],  nodes[702]);
    tranif1 (nodes[558], nodes[324],  nodes[702]);
    tranif1 (nodes[1466], nodes[558],  nodes[702]);
    tranif1 (nodes[558], nodes[546],  nodes[702]);
    tranif1 (nodes[558], nodes[1324],  nodes[702]);
    tranif1 (nodes[558], nodes[179],  nodes[702]);
    tranif1 (nodes[558], nodes[1396],  nodes[702]);
    tranif1 (nodes[558], nodes[167],  nodes[702]);
    tranif1 (nodes[558], nodes[1074],  nodes[702]);
    tranif1 (nodes[558], nodes[1246],  nodes[702]);
    tranif1 (nodes[558], nodes[53],  nodes[702]);
    tranif1 (nodes[558], nodes[691],  nodes[702]);
    tranif1 (nodes[558], nodes[1665],  nodes[702]);
    tranif1 (nodes[191], nodes[558],  nodes[248]);
    tranif1 (nodes[1275], nodes[558],  nodes[778]);
    tranif1 (nodes[558], nodes[687],  nodes[31]);
    tranif1 (nodes[42], nodes[657],  nodes[444]);
    tranif1 (nodes[558], nodes[1196],  nodes[1228]);
    tranif1 (nodes[657], nodes[148],  nodes[1140]);
    tranif1 (nodes[1036], nodes[67],  nodes[943]);
    tranif1 (nodes[558], nodes[1236],  nodes[1632]);
    tranif1 (nodes[558], nodes[1220],  nodes[1632]);
    tranif1 (nodes[558], nodes[1498],  nodes[163]);
    tranif1 (nodes[558], nodes[903],  nodes[163]);
    tranif1 (nodes[558], nodes[1576],  nodes[1620]);
    tranif1 (nodes[862], nodes[1011],  nodes[943]);
    tranif1 (nodes[222], nodes[1687],  nodes[710]);
    tranif1 (nodes[1625], nodes[299],  nodes[710]);
    tranif1 (nodes[169], nodes[1008],  nodes[943]);
    tranif1 (nodes[558], nodes[1714],  nodes[1321]);
    tranif1 (nodes[558], nodes[1103],  nodes[1244]);
    tranif1 (nodes[558], nodes[620],  nodes[1433]);
    tranif1 (nodes[1353], nodes[254],  nodes[710]);
    tranif1 (nodes[1283], nodes[340],  nodes[943]);
    tranif1 (nodes[1023], nodes[433],  nodes[681]);
    tranif1 (nodes[206], nodes[430],  nodes[1446]);
    tranif1 (nodes[558], nodes[311],  nodes[1010]);
    tranif1 (nodes[558], nodes[1334],  nodes[1010]);
    tranif1 (nodes[534], nodes[558],  nodes[1047]);
    tranif1 (nodes[558], nodes[35],  nodes[796]);
    tranif1 (nodes[933], nodes[1407],  nodes[1262]);
    tranif1 (nodes[1490], nodes[296],  nodes[943]);
    tranif1 (nodes[928], nodes[558],  nodes[667]);
    tranif1 (nodes[1032], nodes[891],  nodes[284]);
    tranif1 (nodes[558], nodes[1070],  nodes[292]);
    tranif1 (nodes[558], nodes[60],  nodes[26]);
    tranif1 (nodes[558], nodes[1512],  nodes[26]);
    tranif1 (nodes[558], nodes[1173],  nodes[26]);
    tranif1 (nodes[558], nodes[258],  nodes[26]);
    tranif1 (nodes[558], nodes[245],  nodes[26]);
    tranif1 (nodes[558], nodes[682],  nodes[26]);
    tranif1 (nodes[558], nodes[492],  nodes[26]);
    tranif1 (nodes[558], nodes[1204],  nodes[26]);
    tranif1 (nodes[58], nodes[558],  nodes[26]);
    tranif1 (nodes[558], nodes[342],  nodes[26]);
    tranif1 (nodes[558], nodes[257],  nodes[26]);
    tranif1 (nodes[558], nodes[354],  nodes[26]);
    tranif1 (nodes[558], nodes[1168],  nodes[26]);
    tranif1 (nodes[558], nodes[1721],  nodes[26]);
    tranif1 (nodes[558], nodes[1239],  nodes[26]);
    tranif1 (nodes[461], nodes[558],  nodes[26]);
    tranif1 (nodes[558], nodes[447],  nodes[26]);
    tranif1 (nodes[558], nodes[660],  nodes[26]);
    tranif1 (nodes[558], nodes[1292],  nodes[26]);
    tranif1 (nodes[558], nodes[1114],  nodes[26]);
    tranif1 (nodes[558], nodes[904],  nodes[26]);
    tranif1 (nodes[1419], nodes[558],  nodes[26]);
    tranif1 (nodes[558], nodes[281],  nodes[26]);
    tranif1 (nodes[558], nodes[1164],  nodes[26]);
    tranif1 (nodes[168], nodes[558],  nodes[1651]);
    tranif1 (nodes[704], nodes[1242],  nodes[437]);
    tranif1 (nodes[1104], nodes[889],  nodes[943]);
    tranif1 (nodes[558], nodes[1474],  nodes[991]);
    tranif1 (nodes[558], nodes[48],  nodes[1247]);
    tranif1 (nodes[558], nodes[1331],  nodes[1247]);
    tranif1 (nodes[558], nodes[1039],  nodes[456]);
    tranif1 (nodes[558], nodes[939],  nodes[647]);
    tranif1 (nodes[138], nodes[825],  nodes[943]);
    tranif1 (nodes[558], nodes[717],  nodes[1036]);
    tranif1 (nodes[1650], nodes[558],  nodes[1672]);
    tranif1 (nodes[558], nodes[1270],  nodes[509]);
    tranif1 (nodes[390], nodes[558],  nodes[653]);
    tranif1 (nodes[1455], nodes[558],  nodes[179]);
    tranif1 (nodes[558], nodes[1365],  nodes[862]);
    tranif1 (nodes[9], nodes[657],  nodes[866]);
    tranif1 (nodes[558], nodes[1560],  nodes[1055]);
    tranif1 (nodes[558], nodes[269],  nodes[1038]);
    tranif1 (nodes[1019], nodes[558],  nodes[1622]);
    tranif1 (nodes[558], nodes[1294],  nodes[1622]);
    tranif1 (nodes[1491], nodes[558],  nodes[1484]);
    tranif1 (nodes[1374], nodes[558],  nodes[882]);
    tranif1 (nodes[558], nodes[306],  nodes[725]);
    tranif1 (nodes[558], nodes[1619],  nodes[1448]);
    tranif1 (nodes[858], nodes[831],  nodes[943]);
    tranif1 (nodes[262], nodes[1598],  nodes[1511]);
    tranif1 (nodes[991], nodes[1444],  nodes[1042]);
    tranif1 (nodes[558], nodes[1633],  nodes[172]);
    tranif1 (nodes[657], nodes[210],  nodes[172]);
    tranif1 (nodes[558], nodes[678],  nodes[1357]);
    tranif1 (nodes[1600], nodes[558],  nodes[1302]);
    tranif1 (nodes[1150], nodes[98],  nodes[1186]);
    tranif1 (nodes[964], nodes[558],  nodes[1533]);
    tranif1 (nodes[558], nodes[149],  nodes[331]);
    tranif1 (nodes[1522], nodes[558],  nodes[984]);
    tranif1 (nodes[1399], nodes[558],  nodes[1715]);
    tranif1 (nodes[1399], nodes[558],  nodes[1715]);
    tranif1 (nodes[657], nodes[1105],  nodes[1715]);
    tranif1 (nodes[558], nodes[726],  nodes[677]);
    tranif1 (nodes[558], nodes[565],  nodes[989]);
    tranif1 (nodes[329], nodes[558],  nodes[1022]);
    tranif1 (nodes[1465], nodes[558],  nodes[689]);
    tranif1 (nodes[796], nodes[396],  nodes[943]);
    tranif1 (nodes[1100], nodes[153],  nodes[943]);
    tranif1 (nodes[558], nodes[793],  nodes[1442]);
    tranif1 (nodes[109], nodes[558],  nodes[1380]);
    tranif1 (nodes[405], nodes[558],  nodes[967]);
    tranif1 (nodes[558], nodes[1312],  nodes[1693]);
    tranif1 (nodes[558], nodes[1604],  nodes[1601]);
    tranif1 (nodes[1397], nodes[558],  nodes[1601]);
    tranif1 (nodes[1698], nodes[558],  nodes[1247]);
    tranif1 (nodes[175], nodes[558],  nodes[558]);
    tranif1 (nodes[333], nodes[1030],  nodes[269]);
    tranif1 (nodes[558], nodes[1721],  nodes[603]);
    tranif1 (nodes[336], nodes[1483],  nodes[235]);
    tranif1 (nodes[1084], nodes[558],  nodes[235]);
    tranif1 (nodes[558], nodes[970],  nodes[149]);
    tranif1 (nodes[762], nodes[558],  nodes[149]);
    tranif1 (nodes[478], nodes[558],  nodes[892]);
    tranif1 (nodes[558], nodes[965],  nodes[295]);
    tranif1 (nodes[558], nodes[273],  nodes[791]);
    tranif1 (nodes[558], nodes[677],  nodes[791]);
    tranif1 (nodes[558], nodes[1597],  nodes[116]);
    tranif1 (nodes[1597], nodes[558],  nodes[116]);
    tranif1 (nodes[558], nodes[1597],  nodes[116]);
    tranif1 (nodes[966], nodes[558],  nodes[1683]);
    tranif1 (nodes[558], nodes[325],  nodes[441]);
    tranif1 (nodes[1649], nodes[558],  nodes[1109]);
    tranif1 (nodes[318], nodes[558],  nodes[627]);
    tranif1 (nodes[881], nodes[330],  nodes[538]);
    tranif1 (nodes[1223], nodes[558],  nodes[43]);
    tranif1 (nodes[558], nodes[874],  nodes[282]);
    tranif1 (nodes[1301], nodes[558],  nodes[33]);
    tranif1 (nodes[558], nodes[1517],  nodes[853]);
    tranif1 (nodes[558], nodes[1388],  nodes[425]);
    tranif1 (nodes[558], nodes[295],  nodes[425]);
    tranif1 (nodes[558], nodes[1584],  nodes[876]);
    tranif1 (nodes[833], nodes[1458],  nodes[283]);
    tranif1 (nodes[558], nodes[326],  nodes[1356]);
    tranif1 (nodes[558], nodes[637],  nodes[1318]);
    tranif1 (nodes[558], nodes[516],  nodes[1691]);
    tranif1 (nodes[401], nodes[558],  nodes[394]);
    tranif1 (nodes[471], nodes[558],  nodes[1415]);
    tranif1 (nodes[466], nodes[558],  nodes[1415]);
    tranif1 (nodes[698], nodes[1290],  nodes[710]);
    tranif1 (nodes[955], nodes[111],  nodes[943]);
    tranif1 (nodes[1690], nodes[62],  nodes[943]);
    tranif1 (nodes[1669], nodes[374],  nodes[943]);
    tranif1 (nodes[558], nodes[888],  nodes[675]);
    tranif1 (nodes[558], nodes[888],  nodes[675]);
    tranif1 (nodes[872], nodes[558],  nodes[697]);
    tranif1 (nodes[558], nodes[636],  nodes[1239]);
    tranif1 (nodes[106], nodes[732],  nodes[792]);
    tranif1 (nodes[93], nodes[558],  nodes[1005]);
    tranif1 (nodes[558], nodes[419],  nodes[978]);
    tranif1 (nodes[1320], nodes[558],  nodes[1328]);
    tranif1 (nodes[1688], nodes[558],  nodes[1304]);
    tranif1 (nodes[998], nodes[558],  nodes[828]);
    tranif1 (nodes[558], nodes[1145],  nodes[248]);
    tranif1 (nodes[558], nodes[604],  nodes[248]);
    tranif1 (nodes[599], nodes[533],  nodes[710]);
    tranif1 (nodes[694], nodes[558],  nodes[1064]);
    tranif1 (nodes[849], nodes[558],  nodes[321]);
    tranif1 (nodes[247], nodes[657],  nodes[321]);
    tranif1 (nodes[558], nodes[384],  nodes[1228]);
    tranif1 (nodes[558], nodes[384],  nodes[1228]);
    tranif1 (nodes[558], nodes[385],  nodes[1377]);
    tranif1 (nodes[1614], nodes[558],  nodes[1177]);
    tranif1 (nodes[300], nodes[558],  nodes[857]);
    tranif1 (nodes[520], nodes[558],  nodes[353]);
    tranif1 (nodes[520], nodes[558],  nodes[353]);
    tranif1 (nodes[224], nodes[558],  nodes[353]);
    tranif1 (nodes[558], nodes[60],  nodes[194]);
    tranif1 (nodes[558], nodes[1512],  nodes[194]);
    tranif1 (nodes[558], nodes[84],  nodes[194]);
    tranif1 (nodes[1623], nodes[558],  nodes[194]);
    tranif1 (nodes[403], nodes[558],  nodes[194]);
    tranif1 (nodes[1428], nodes[558],  nodes[194]);
    tranif1 (nodes[492], nodes[558],  nodes[194]);
    tranif1 (nodes[1204], nodes[558],  nodes[194]);
    tranif1 (nodes[558], nodes[1259],  nodes[194]);
    tranif1 (nodes[342], nodes[558],  nodes[194]);
    tranif1 (nodes[1355], nodes[558],  nodes[194]);
    tranif1 (nodes[787], nodes[558],  nodes[194]);
    tranif1 (nodes[575], nodes[558],  nodes[194]);
    tranif1 (nodes[558], nodes[1243],  nodes[194]);
    tranif1 (nodes[558], nodes[822],  nodes[194]);
    tranif1 (nodes[558], nodes[1420],  nodes[194]);
    tranif1 (nodes[1342], nodes[558],  nodes[194]);
    tranif1 (nodes[1504], nodes[558],  nodes[194]);
    tranif1 (nodes[558], nodes[1168],  nodes[194]);
    tranif1 (nodes[558], nodes[145],  nodes[194]);
    tranif1 (nodes[558], nodes[1524],  nodes[194]);
    tranif1 (nodes[558], nodes[1210],  nodes[194]);
    tranif1 (nodes[558], nodes[461],  nodes[194]);
    tranif1 (nodes[1155], nodes[558],  nodes[194]);
    tranif1 (nodes[301], nodes[558],  nodes[194]);
    tranif1 (nodes[1385], nodes[558],  nodes[194]);
    tranif1 (nodes[650], nodes[558],  nodes[558]);
    tranif1 (nodes[944], nodes[558],  nodes[759]);
    tranif1 (nodes[343], nodes[1300],  nodes[879]);
    tranif1 (nodes[664], nodes[558],  nodes[1006]);
    tranif1 (nodes[330], nodes[675],  nodes[710]);
    tranif1 (nodes[558], nodes[612],  nodes[353]);
    tranif1 (nodes[558], nodes[612],  nodes[353]);
    tranif1 (nodes[294], nodes[14],  nodes[943]);
    tranif1 (nodes[832], nodes[586],  nodes[943]);
    tranif1 (nodes[60], nodes[558],  nodes[1567]);
    tranif1 (nodes[1487], nodes[558],  nodes[1567]);
    tranif1 (nodes[1031], nodes[558],  nodes[1567]);
    tranif1 (nodes[558], nodes[1428],  nodes[1567]);
    tranif1 (nodes[58], nodes[558],  nodes[1567]);
    tranif1 (nodes[342], nodes[558],  nodes[1567]);
    tranif1 (nodes[558], nodes[1381],  nodes[1567]);
    tranif1 (nodes[579], nodes[558],  nodes[1567]);
    tranif1 (nodes[120], nodes[558],  nodes[1567]);
    tranif1 (nodes[677], nodes[558],  nodes[1567]);
    tranif1 (nodes[447], nodes[558],  nodes[1567]);
    tranif1 (nodes[660], nodes[558],  nodes[1567]);
    tranif1 (nodes[1430], nodes[558],  nodes[1567]);
    tranif1 (nodes[558], nodes[904],  nodes[1567]);
    tranif1 (nodes[607], nodes[558],  nodes[1567]);
    tranif1 (nodes[150], nodes[613],  nodes[1682]);
    tranif1 (nodes[1256], nodes[558],  nodes[91]);
    tranif1 (nodes[574], nodes[657],  nodes[91]);
    tranif1 (nodes[543], nodes[558],  nodes[339]);
    tranif1 (nodes[558], nodes[239],  nodes[595]);
    tranif1 (nodes[558], nodes[992],  nodes[595]);
    tranif1 (nodes[859], nodes[558],  nodes[1247]);
    tranif1 (nodes[907], nodes[676],  nodes[943]);
    tranif1 (nodes[1536], nodes[657],  nodes[17]);
    tranif1 (nodes[646], nodes[558],  nodes[17]);
    tranif1 (nodes[889], nodes[558],  nodes[1114]);
    tranif1 (nodes[558], nodes[327],  nodes[1226]);
    tranif1 (nodes[1661], nodes[684],  nodes[1564]);
    tranif1 (nodes[1095], nodes[1437],  nodes[1564]);
    tranif1 (nodes[87], nodes[1282],  nodes[1564]);
    tranif1 (nodes[1424], nodes[1242],  nodes[1564]);
    tranif1 (nodes[719], nodes[413],  nodes[1564]);
    tranif1 (nodes[558], nodes[1322],  nodes[320]);
    tranif1 (nodes[558], nodes[735],  nodes[320]);
    tranif1 (nodes[471], nodes[558],  nodes[353]);
    tranif1 (nodes[471], nodes[558],  nodes[353]);
    tranif1 (nodes[595], nodes[558],  nodes[354]);
    tranif1 (nodes[558], nodes[643],  nodes[444]);
    tranif1 (nodes[558], nodes[1613],  nodes[444]);
    tranif1 (nodes[1134], nodes[1431],  nodes[943]);
    tranif1 (nodes[256], nodes[558],  nodes[1478]);
    tranif1 (nodes[558], nodes[924],  nodes[1313]);
    tranif1 (nodes[710], nodes[558],  nodes[1105]);
    tranif1 (nodes[710], nodes[558],  nodes[1105]);
    tranif1 (nodes[558], nodes[710],  nodes[1105]);
    tranif1 (nodes[710], nodes[558],  nodes[1105]);
    tranif1 (nodes[558], nodes[710],  nodes[1105]);
    tranif1 (nodes[545], nodes[558],  nodes[1488]);
    tranif1 (nodes[1547], nodes[558],  nodes[1488]);
    tranif1 (nodes[815], nodes[558],  nodes[45]);
    tranif1 (nodes[570], nodes[558],  nodes[647]);
    tranif1 (nodes[1287], nodes[1491],  nodes[801]);
    tranif1 (nodes[558], nodes[467],  nodes[470]);
    tranif1 (nodes[737], nodes[146],  nodes[943]);
    tranif1 (nodes[1531], nodes[1188],  nodes[801]);
    tranif1 (nodes[558], nodes[513],  nodes[885]);
    tranif1 (nodes[37], nodes[558],  nodes[353]);
    tranif1 (nodes[37], nodes[558],  nodes[353]);
    tranif1 (nodes[313], nodes[350],  nodes[96]);
    tranif1 (nodes[558], nodes[649],  nodes[96]);
    tranif1 (nodes[798], nodes[558],  nodes[288]);
    tranif1 (nodes[794], nodes[657],  nodes[288]);
    tranif1 (nodes[657], nodes[826],  nodes[1429]);
    tranif1 (nodes[558], nodes[625],  nodes[43]);
    tranif1 (nodes[34], nodes[558],  nodes[1532]);
    tranif1 (nodes[652], nodes[558],  nodes[751]);
    tranif1 (nodes[475], nodes[558],  nodes[1677]);
    tranif1 (nodes[999], nodes[657],  nodes[1677]);
    tranif1 (nodes[958], nodes[865],  nodes[943]);
    tranif1 (nodes[85], nodes[1405],  nodes[1186]);
    tranif1 (nodes[1188], nodes[1648],  nodes[1186]);
    tranif1 (nodes[1287], nodes[1],  nodes[1186]);
    tranif1 (nodes[1067], nodes[558],  nodes[582]);
    tranif1 (nodes[657], nodes[821],  nodes[582]);
    tranif1 (nodes[448], nodes[1336],  nodes[1186]);
    tranif1 (nodes[166], nodes[589],  nodes[1186]);
    tranif1 (nodes[263], nodes[558],  nodes[1629]);
    tranif1 (nodes[1502], nodes[558],  nodes[707]);
    tranif1 (nodes[654], nodes[558],  nodes[71]);
    tranif1 (nodes[1001], nodes[777],  nodes[1186]);
    tranif1 (nodes[558], nodes[1719],  nodes[858]);
    tranif1 (nodes[558], nodes[1717],  nodes[60]);
    tranif1 (nodes[945], nodes[657],  nodes[520]);
    tranif1 (nodes[945], nodes[657],  nodes[520]);
    tranif1 (nodes[558], nodes[253],  nodes[1104]);
    tranif1 (nodes[558], nodes[362],  nodes[1552]);
    tranif1 (nodes[558], nodes[797],  nodes[892]);
    tranif1 (nodes[558], nodes[678],  nodes[644]);
    tranif1 (nodes[558], nodes[854],  nodes[975]);
    tranif1 (nodes[803], nodes[558],  nodes[1084]);
    tranif1 (nodes[558], nodes[1314],  nodes[1084]);
    tranif1 (nodes[1494], nodes[1454],  nodes[1205]);
    tranif1 (nodes[558], nodes[260],  nodes[1205]);
    tranif1 (nodes[982], nodes[1689],  nodes[943]);
    tranif1 (nodes[657], nodes[1001],  nodes[943]);
    tranif1 (nodes[88], nodes[522],  nodes[943]);
    tranif1 (nodes[914], nodes[484],  nodes[1386]);
    tranif1 (nodes[558], nodes[307],  nodes[31]);
    tranif1 (nodes[558], nodes[1580],  nodes[1287]);
    tranif1 (nodes[558], nodes[1580],  nodes[1287]);
    tranif1 (nodes[558], nodes[435],  nodes[86]);
    tranif1 (nodes[435], nodes[558],  nodes[86]);
    tranif1 (nodes[435], nodes[558],  nodes[86]);
    tranif1 (nodes[435], nodes[558],  nodes[86]);
    tranif1 (nodes[248], nodes[1624],  nodes[710]);
    tranif1 (nodes[558], nodes[616],  nodes[286]);
    tranif1 (nodes[558], nodes[482],  nodes[803]);
    tranif1 (nodes[736], nodes[558],  nodes[210]);
    tranif1 (nodes[736], nodes[558],  nodes[210]);
    tranif1 (nodes[736], nodes[558],  nodes[210]);
    tranif1 (nodes[736], nodes[558],  nodes[210]);
    tranif1 (nodes[558], nodes[959],  nodes[294]);
    tranif1 (nodes[1592], nodes[558],  nodes[128]);
    tranif1 (nodes[42], nodes[558],  nodes[353]);
    tranif1 (nodes[42], nodes[558],  nodes[353]);
    tranif1 (nodes[1613], nodes[558],  nodes[353]);
    tranif1 (nodes[1165], nodes[558],  nodes[910]);
    tranif1 (nodes[989], nodes[658],  nodes[943]);
    tranif1 (nodes[558], nodes[1304],  nodes[673]);
    tranif1 (nodes[558], nodes[39],  nodes[15]);
    tranif1 (nodes[880], nodes[1514],  nodes[710]);
    tranif1 (nodes[558], nodes[549],  nodes[708]);
    tranif1 (nodes[1531], nodes[305],  nodes[943]);
    tranif1 (nodes[629], nodes[202],  nodes[480]);
    tranif1 (nodes[1606], nodes[472],  nodes[710]);
    tranif1 (nodes[90], nodes[44],  nodes[943]);
    tranif1 (nodes[229], nodes[558],  nodes[683]);
    tranif1 (nodes[558], nodes[1380],  nodes[1154]);
    tranif1 (nodes[347], nodes[558],  nodes[904]);
    tranif1 (nodes[608], nodes[559],  nodes[943]);
    tranif1 (nodes[373], nodes[558],  nodes[353]);
    tranif1 (nodes[373], nodes[558],  nodes[353]);
    tranif1 (nodes[1720], nodes[558],  nodes[353]);
    tranif1 (nodes[657], nodes[54],  nodes[943]);
    tranif1 (nodes[68], nodes[722],  nodes[943]);
    tranif1 (nodes[302], nodes[558],  nodes[409]);
    tranif1 (nodes[957], nodes[841],  nodes[362]);
    tranif1 (nodes[681], nodes[250],  nodes[362]);
    tranif1 (nodes[740], nodes[350],  nodes[362]);
    tranif1 (nodes[1063], nodes[1071],  nodes[362]);
    tranif1 (nodes[477], nodes[296],  nodes[362]);
    tranif1 (nodes[336], nodes[277],  nodes[362]);
    tranif1 (nodes[1318], nodes[722],  nodes[362]);
    tranif1 (nodes[875], nodes[469],  nodes[943]);
    tranif1 (nodes[558], nodes[844],  nodes[1664]);
    tranif1 (nodes[1287], nodes[573],  nodes[325]);
    tranif1 (nodes[450], nodes[1656],  nodes[613]);
    tranif1 (nodes[1159], nodes[558],  nodes[613]);
    tranif1 (nodes[493], nodes[657],  nodes[943]);
    tranif1 (nodes[1452], nodes[1481],  nodes[943]);
    tranif1 (nodes[808], nodes[560],  nodes[943]);
    tranif1 (nodes[558], nodes[1517],  nodes[572]);
    tranif1 (nodes[1525], nodes[1348],  nodes[693]);
    tranif1 (nodes[558], nodes[169],  nodes[139]);
    tranif1 (nodes[1421], nodes[558],  nodes[334]);
    tranif1 (nodes[558], nodes[643],  nodes[353]);
    tranif1 (nodes[558], nodes[643],  nodes[353]);
    tranif1 (nodes[558], nodes[46],  nodes[248]);
    tranif1 (nodes[1185], nodes[558],  nodes[1137]);
    tranif1 (nodes[412], nodes[558],  nodes[560]);
    tranif1 (nodes[558], nodes[274],  nodes[860]);
    tranif1 (nodes[85], nodes[436],  nodes[943]);
    tranif1 (nodes[1284], nodes[896],  nodes[943]);
    tranif1 (nodes[180], nodes[558],  nodes[1716]);
    tranif1 (nodes[558], nodes[588],  nodes[1349]);
    tranif1 (nodes[1370], nodes[558],  nodes[1045]);
    tranif1 (nodes[132], nodes[1321],  nodes[943]);
    tranif1 (nodes[1307], nodes[1254],  nodes[943]);
    tranif1 (nodes[558], nodes[1347],  nodes[550]);
    tranif1 (nodes[816], nodes[1137],  nodes[790]);
    tranif1 (nodes[697], nodes[250],  nodes[943]);
    tranif1 (nodes[864], nodes[825],  nodes[639]);
    tranif1 (nodes[1588], nodes[558],  nodes[175]);
    tranif1 (nodes[1417], nodes[558],  nodes[747]);
    tranif1 (nodes[1309], nodes[558],  nodes[1460]);
    tranif1 (nodes[558], nodes[201],  nodes[1174]);
    tranif1 (nodes[798], nodes[558],  nodes[353]);
    tranif1 (nodes[798], nodes[558],  nodes[353]);
    tranif1 (nodes[288], nodes[558],  nodes[353]);
    tranif1 (nodes[525], nodes[558],  nodes[943]);
    tranif1 (nodes[628], nodes[558],  nodes[943]);
    tranif1 (nodes[558], nodes[1470],  nodes[1111]);
    tranif1 (nodes[1614], nodes[558],  nodes[1111]);
    tranif1 (nodes[558], nodes[313],  nodes[1680]);
    tranif1 (nodes[558], nodes[649],  nodes[1680]);
    tranif1 (nodes[558], nodes[984],  nodes[956]);
    tranif1 (nodes[242], nodes[558],  nodes[1521]);
    tranif1 (nodes[1150], nodes[1148],  nodes[325]);
    tranif1 (nodes[504], nodes[137],  nodes[440]);
    tranif1 (nodes[558], nodes[1649],  nodes[1382]);
    tranif1 (nodes[558], nodes[300],  nodes[1382]);
    tranif1 (nodes[558], nodes[1433],  nodes[90]);
    tranif1 (nodes[256], nodes[558],  nodes[120]);
    tranif1 (nodes[185], nodes[1063],  nodes[1645]);
    tranif1 (nodes[558], nodes[404],  nodes[1645]);
    tranif1 (nodes[1352], nodes[558],  nodes[1258]);
    tranif1 (nodes[1169], nodes[558],  nodes[987]);
    tranif1 (nodes[531], nodes[558],  nodes[95]);
    tranif1 (nodes[1051], nodes[31],  nodes[943]);
    tranif1 (nodes[1149], nodes[1368],  nodes[710]);
    tranif1 (nodes[558], nodes[612],  nodes[1453]);
    tranif1 (nodes[558], nodes[1720],  nodes[1453]);
    tranif1 (nodes[113], nodes[558],  nodes[126]);
    tranif1 (nodes[558], nodes[1391],  nodes[750]);
    tranif1 (nodes[1610], nodes[558],  nodes[640]);
    tranif1 (nodes[532], nodes[558],  nodes[1217]);
    tranif1 (nodes[558], nodes[476],  nodes[43]);
    tranif1 (nodes[1213], nodes[558],  nodes[453]);
    tranif1 (nodes[558], nodes[620],  nodes[1371]);
    tranif1 (nodes[558], nodes[51],  nodes[439]);
    tranif1 (nodes[334], nodes[558],  nodes[1553]);
    tranif1 (nodes[605], nodes[558],  nodes[1002]);
    tranif1 (nodes[605], nodes[558],  nodes[1002]);
    tranif1 (nodes[558], nodes[1541],  nodes[1477]);
    tranif1 (nodes[1107], nodes[558],  nodes[1428]);
    tranif1 (nodes[604], nodes[558],  nodes[1428]);
    tranif1 (nodes[89], nodes[558],  nodes[558]);
    tranif1 (nodes[272], nodes[558],  nodes[646]);
    tranif1 (nodes[1293], nodes[558],  nodes[1174]);
    tranif1 (nodes[1455], nodes[558],  nodes[131]);
    tranif1 (nodes[558], nodes[1331],  nodes[800]);
    tranif1 (nodes[741], nodes[558],  nodes[1247]);
    tranif1 (nodes[1014], nodes[121],  nodes[1564]);
    tranif1 (nodes[1387], nodes[1630],  nodes[1564]);
    tranif1 (nodes[266], nodes[1037],  nodes[943]);
    tranif1 (nodes[650], nodes[657],  nodes[42]);
    tranif1 (nodes[650], nodes[657],  nodes[42]);
    tranif1 (nodes[973], nodes[558],  nodes[1702]);
    tranif1 (nodes[1119], nodes[558],  nodes[1471]);
    tranif1 (nodes[621], nodes[1586],  nodes[943]);
    tranif1 (nodes[1046], nodes[577],  nodes[710]);
    tranif1 (nodes[956], nodes[558],  nodes[476]);
    tranif1 (nodes[657], nodes[984],  nodes[476]);
    tranif1 (nodes[558], nodes[1244],  nodes[1562]);
    tranif1 (nodes[558], nodes[1351],  nodes[1562]);
    tranif1 (nodes[558], nodes[961],  nodes[1503]);
    tranif1 (nodes[226], nodes[1093],  nodes[710]);
    tranif1 (nodes[558], nodes[1358],  nodes[245]);
    tranif1 (nodes[558], nodes[14],  nodes[671]);
    tranif1 (nodes[1662], nodes[558],  nodes[1124]);
    tranif1 (nodes[1401], nodes[558],  nodes[1269]);
    tranif1 (nodes[1249], nodes[558],  nodes[1269]);
    tranif1 (nodes[1451], nodes[668],  nodes[821]);
    tranif1 (nodes[558], nodes[1593],  nodes[226]);
    tranif1 (nodes[558], nodes[196],  nodes[543]);
    tranif1 (nodes[1468], nodes[657],  nodes[543]);
    tranif1 (nodes[236], nodes[558],  nodes[1708]);
    tranif1 (nodes[657], nodes[1237],  nodes[475]);
    tranif1 (nodes[558], nodes[827],  nodes[1350]);
    tranif1 (nodes[1472], nodes[827],  nodes[710]);
    tranif1 (nodes[1581], nodes[1275],  nodes[710]);
    tranif1 (nodes[1133], nodes[558],  nodes[1626]);
    tranif1 (nodes[702], nodes[558],  nodes[1626]);
    tranif1 (nodes[1353], nodes[1128],  nodes[821]);
    tranif1 (nodes[1037], nodes[558],  nodes[1086]);
    tranif1 (nodes[1105], nodes[558],  nodes[1399]);
    tranif1 (nodes[972], nodes[558],  nodes[319]);
    tranif1 (nodes[425], nodes[558],  nodes[936]);
    tranif1 (nodes[1005], nodes[657],  nodes[1325]);
    tranif1 (nodes[657], nodes[1005],  nodes[1325]);
    tranif1 (nodes[611], nodes[558],  nodes[43]);
    tranif1 (nodes[1106], nodes[558],  nodes[245]);
    tranif1 (nodes[1350], nodes[50],  nodes[710]);
    tranif1 (nodes[558], nodes[36],  nodes[600]);
    tranif1 (nodes[1048], nodes[558],  nodes[1721]);
    tranif1 (nodes[935], nodes[1636],  nodes[710]);
    tranif1 (nodes[558], nodes[503],  nodes[1394]);
    tranif1 (nodes[280], nodes[1630],  nodes[1468]);
    tranif1 (nodes[3], nodes[1437],  nodes[1468]);
    tranif1 (nodes[998], nodes[684],  nodes[1468]);
    tranif1 (nodes[1389], nodes[1242],  nodes[1468]);
    tranif1 (nodes[558], nodes[1004],  nodes[1408]);
    tranif1 (nodes[558], nodes[553],  nodes[1662]);
    tranif1 (nodes[1299], nodes[721],  nodes[1468]);
    tranif1 (nodes[558], nodes[1347],  nodes[862]);
    tranif1 (nodes[376], nodes[558],  nodes[107]);
    tranif1 (nodes[1151], nodes[182],  nodes[236]);
    tranif1 (nodes[141], nodes[558],  nodes[124]);
    tranif1 (nodes[1215], nodes[1528],  nodes[710]);
    tranif1 (nodes[109], nodes[1161],  nodes[710]);
    tranif1 (nodes[1198], nodes[626],  nodes[1401]);
    tranif1 (nodes[391], nodes[558],  nodes[529]);
    tranif1 (nodes[391], nodes[558],  nodes[529]);
    tranif1 (nodes[391], nodes[558],  nodes[529]);
    tranif1 (nodes[19], nodes[558],  nodes[770]);
    tranif1 (nodes[657], nodes[1150],  nodes[943]);
    tranif1 (nodes[265], nodes[182],  nodes[943]);
    tranif1 (nodes[1211], nodes[897],  nodes[943]);
    tranif1 (nodes[558], nodes[368],  nodes[446]);
    tranif1 (nodes[1354], nodes[558],  nodes[1165]);
    tranif1 (nodes[879], nodes[558],  nodes[1214]);
    tranif1 (nodes[558], nodes[1635],  nodes[966]);
    tranif1 (nodes[203], nodes[657],  nodes[966]);
    tranif1 (nodes[558], nodes[770],  nodes[559]);
    tranif1 (nodes[558], nodes[1271],  nodes[1596]);
    tranif1 (nodes[140], nodes[657],  nodes[1596]);
    tranif1 (nodes[1242], nodes[657],  nodes[943]);
    tranif1 (nodes[114], nodes[1402],  nodes[943]);
    tranif1 (nodes[1116], nodes[1014],  nodes[710]);
    tranif1 (nodes[1495], nodes[1546],  nodes[1600]);
    tranif1 (nodes[558], nodes[1044],  nodes[31]);
    tranif1 (nodes[979], nodes[558],  nodes[905]);
    tranif1 (nodes[558], nodes[156],  nodes[1533]);
    tranif1 (nodes[175], nodes[657],  nodes[373]);
    tranif1 (nodes[175], nodes[657],  nodes[373]);
    tranif1 (nodes[267], nodes[558],  nodes[1175]);
    tranif1 (nodes[657], nodes[1473],  nodes[943]);
    tranif1 (nodes[558], nodes[882],  nodes[597]);
    tranif1 (nodes[558], nodes[1056],  nodes[761]);
    tranif1 (nodes[619], nodes[695],  nodes[78]);
    tranif1 (nodes[1179], nodes[558],  nodes[78]);
    tranif1 (nodes[745], nodes[674],  nodes[943]);
    tranif1 (nodes[512], nodes[1130],  nodes[943]);
    tranif1 (nodes[1099], nodes[1102],  nodes[943]);
    tranif1 (nodes[558], nodes[269],  nodes[1241]);
    tranif1 (nodes[298], nodes[558],  nodes[353]);
    tranif1 (nodes[298], nodes[558],  nodes[353]);
    tranif1 (nodes[23], nodes[558],  nodes[353]);
    tranif1 (nodes[558], nodes[1279],  nodes[600]);
    tranif1 (nodes[969], nodes[558],  nodes[161]);
    tranif1 (nodes[801], nodes[657],  nodes[161]);
    tranif1 (nodes[558], nodes[715],  nodes[641]);
    tranif1 (nodes[558], nodes[1704],  nodes[641]);
    tranif1 (nodes[654], nodes[558],  nodes[1247]);
    tranif1 (nodes[604], nodes[558],  nodes[804]);
    tranif1 (nodes[166], nodes[615],  nodes[325]);
    tranif1 (nodes[1042], nodes[558],  nodes[1577]);
    tranif1 (nodes[414], nodes[558],  nodes[1043]);
    tranif1 (nodes[1001], nodes[843],  nodes[325]);
    tranif1 (nodes[558], nodes[1257],  nodes[1218]);
    tranif1 (nodes[558], nodes[1587],  nodes[894]);
    tranif1 (nodes[490], nodes[558],  nodes[1393]);
    tranif1 (nodes[557], nodes[1073],  nodes[344]);
    tranif1 (nodes[230], nodes[657],  nodes[826]);
    tranif1 (nodes[585], nodes[20],  nodes[344]);
    tranif1 (nodes[1316], nodes[558],  nodes[344]);
    tranif1 (nodes[934], nodes[73],  nodes[943]);
    tranif1 (nodes[558], nodes[1465],  nodes[248]);
    tranif1 (nodes[558], nodes[1349],  nodes[1501]);
    tranif1 (nodes[558], nodes[1349],  nodes[1501]);
    tranif1 (nodes[1349], nodes[558],  nodes[1501]);
    tranif1 (nodes[558], nodes[1349],  nodes[1501]);
    tranif1 (nodes[160], nodes[1049],  nodes[943]);
    tranif1 (nodes[558], nodes[647],  nodes[477]);
    tranif1 (nodes[264], nodes[558],  nodes[1149]);
    tranif1 (nodes[1218], nodes[558],  nodes[1565]);
    tranif1 (nodes[1218], nodes[558],  nodes[1565]);
    tranif1 (nodes[1276], nodes[248],  nodes[710]);
    tranif1 (nodes[501], nodes[1713],  nodes[943]);
    tranif1 (nodes[558], nodes[1512],  nodes[971]);
    tranif1 (nodes[558], nodes[258],  nodes[971]);
    tranif1 (nodes[558], nodes[84],  nodes[971]);
    tranif1 (nodes[558], nodes[788],  nodes[971]);
    tranif1 (nodes[558], nodes[1057],  nodes[971]);
    tranif1 (nodes[558], nodes[204],  nodes[971]);
    tranif1 (nodes[558], nodes[1582],  nodes[971]);
    tranif1 (nodes[558], nodes[1204],  nodes[971]);
    tranif1 (nodes[558], nodes[712],  nodes[971]);
    tranif1 (nodes[558], nodes[157],  nodes[971]);
    tranif1 (nodes[558], nodes[1086],  nodes[971]);
    tranif1 (nodes[558], nodes[487],  nodes[971]);
    tranif1 (nodes[558], nodes[1239],  nodes[971]);
    tranif1 (nodes[558], nodes[285],  nodes[971]);
    tranif1 (nodes[558], nodes[1524],  nodes[971]);
    tranif1 (nodes[558], nodes[273],  nodes[971]);
    tranif1 (nodes[558], nodes[750],  nodes[971]);
    tranif1 (nodes[558], nodes[932],  nodes[971]);
    tranif1 (nodes[558], nodes[309],  nodes[971]);
    tranif1 (nodes[558], nodes[219],  nodes[971]);
    tranif1 (nodes[1091], nodes[1360],  nodes[710]);
    tranif1 (nodes[1106], nodes[558],  nodes[84]);
    tranif1 (nodes[1262], nodes[558],  nodes[1679]);
    tranif1 (nodes[504], nodes[1438],  nodes[943]);
    tranif1 (nodes[1574], nodes[1228],  nodes[943]);
    tranif1 (nodes[1640], nodes[558],  nodes[843]);
    tranif1 (nodes[702], nodes[119],  nodes[943]);
    tranif1 (nodes[558], nodes[1006],  nodes[328]);
    tranif1 (nodes[119], nodes[237],  nodes[879]);
    tranif1 (nodes[310], nodes[724],  nodes[879]);
    tranif1 (nodes[1272], nodes[248],  nodes[710]);
    tranif1 (nodes[270], nodes[558],  nodes[503]);
    tranif1 (nodes[558], nodes[1684],  nodes[833]);
    tranif1 (nodes[256], nodes[558],  nodes[0]);
    tranif1 (nodes[1303], nodes[508],  nodes[335]);
    tranif1 (nodes[558], nodes[1460],  nodes[1669]);
    tranif1 (nodes[452], nodes[681],  nodes[704]);
    tranif1 (nodes[558], nodes[1691],  nodes[704]);
    tranif1 (nodes[737], nodes[54],  nodes[534]);
    tranif1 (nodes[1234], nodes[1009],  nodes[534]);
    tranif1 (nodes[450], nodes[978],  nodes[534]);
    tranif1 (nodes[162], nodes[1475],  nodes[534]);
    tranif1 (nodes[727], nodes[1405],  nodes[534]);
    tranif1 (nodes[858], nodes[263],  nodes[534]);
    tranif1 (nodes[1136], nodes[679],  nodes[534]);
    tranif1 (nodes[1653], nodes[1494],  nodes[534]);
    tranif1 (nodes[1028], nodes[558],  nodes[251]);
    tranif1 (nodes[558], nodes[353],  nodes[251]);
    tranif1 (nodes[558], nodes[353],  nodes[251]);
    tranif1 (nodes[353], nodes[558],  nodes[251]);
    tranif1 (nodes[353], nodes[558],  nodes[251]);
    tranif1 (nodes[558], nodes[19],  nodes[1708]);
    tranif1 (nodes[1108], nodes[54],  nodes[1060]);
    tranif1 (nodes[991], nodes[1150],  nodes[1060]);
    tranif1 (nodes[1287], nodes[1473],  nodes[1060]);
    tranif1 (nodes[1302], nodes[1188],  nodes[1060]);
    tranif1 (nodes[1405], nodes[892],  nodes[1060]);
    tranif1 (nodes[166], nodes[1503],  nodes[1060]);
    tranif1 (nodes[1336], nodes[833],  nodes[1060]);
    tranif1 (nodes[493], nodes[1001],  nodes[1060]);
    tranif1 (nodes[1124], nodes[1065],  nodes[943]);
    tranif1 (nodes[558], nodes[1144],  nodes[1571]);
    tranif1 (nodes[439], nodes[558],  nodes[1194]);
    tranif1 (nodes[1178], nodes[558],  nodes[848]);
    tranif1 (nodes[398], nodes[824],  nodes[943]);
    tranif1 (nodes[558], nodes[728],  nodes[1465]);
    tranif1 (nodes[1372], nodes[972],  nodes[388]);
    tranif1 (nodes[1250], nodes[558],  nodes[825]);
    tranif1 (nodes[742], nodes[558],  nodes[943]);
    tranif1 (nodes[454], nodes[558],  nodes[616]);
    tranif1 (nodes[774], nodes[558],  nodes[1419]);
    tranif1 (nodes[558], nodes[1258],  nodes[390]);
    tranif1 (nodes[558], nodes[1415],  nodes[1418]);
    tranif1 (nodes[1299], nodes[1147],  nodes[1564]);
    tranif1 (nodes[922], nodes[558],  nodes[620]);
    tranif1 (nodes[558], nodes[1115],  nodes[620]);
    tranif1 (nodes[1238], nodes[558],  nodes[1295]);
    tranif1 (nodes[1060], nodes[657],  nodes[1295]);
    tranif1 (nodes[663], nodes[1209],  nodes[943]);
    tranif1 (nodes[69], nodes[1181],  nodes[710]);
    tranif1 (nodes[171], nodes[28],  nodes[943]);
    tranif1 (nodes[558], nodes[437],  nodes[1247]);
    tranif1 (nodes[558], nodes[252],  nodes[1710]);
    tranif1 (nodes[558], nodes[1339],  nodes[799]);
    tranif1 (nodes[650], nodes[558],  nodes[643]);
    tranif1 (nodes[650], nodes[558],  nodes[643]);
    tranif1 (nodes[650], nodes[558],  nodes[643]);
    tranif1 (nodes[558], nodes[650],  nodes[643]);
    tranif1 (nodes[558], nodes[650],  nodes[643]);
    tranif1 (nodes[650], nodes[558],  nodes[643]);
    tranif1 (nodes[650], nodes[558],  nodes[643]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[1156], nodes[657],  nodes[102]);
    tranif1 (nodes[592], nodes[558],  nodes[1314]);
    tranif1 (nodes[1617], nodes[1327],  nodes[1314]);
    tranif1 (nodes[558], nodes[302],  nodes[1083]);
    tranif1 (nodes[558], nodes[1019],  nodes[1083]);
    tranif1 (nodes[648], nodes[558],  nodes[1200]);
    tranif1 (nodes[558], nodes[548],  nodes[1435]);
    tranif1 (nodes[558], nodes[1277],  nodes[1020]);
    tranif1 (nodes[558], nodes[1723],  nodes[1436]);
    tranif1 (nodes[1614], nodes[558],  nodes[1436]);
    tranif1 (nodes[903], nodes[1631],  nodes[1184]);
    tranif1 (nodes[657], nodes[1651],  nodes[943]);
    tranif1 (nodes[1172], nodes[1085],  nodes[372]);
    tranif1 (nodes[1290], nodes[912],  nodes[248]);
    tranif1 (nodes[773], nodes[558],  nodes[273]);
    tranif1 (nodes[17], nodes[558],  nodes[964]);
    tranif1 (nodes[1536], nodes[558],  nodes[964]);
    tranif1 (nodes[535], nodes[558],  nodes[663]);
    tranif1 (nodes[558], nodes[1286],  nodes[470]);
    tranif1 (nodes[558], nodes[135],  nodes[127]);
    tranif1 (nodes[901], nodes[558],  nodes[872]);
    tranif1 (nodes[1723], nodes[299],  nodes[1245]);
    tranif1 (nodes[657], nodes[1340],  nodes[1152]);
    tranif1 (nodes[657], nodes[1340],  nodes[1152]);
    tranif1 (nodes[1340], nodes[657],  nodes[1152]);
    tranif1 (nodes[1340], nodes[657],  nodes[1152]);
    tranif1 (nodes[657], nodes[1340],  nodes[1152]);
    tranif1 (nodes[558], nodes[1081],  nodes[1560]);
    tranif1 (nodes[558], nodes[1329],  nodes[1609]);
    tranif1 (nodes[558], nodes[1499],  nodes[1450]);
    tranif1 (nodes[1712], nodes[558],  nodes[926]);
    tranif1 (nodes[566], nodes[661],  nodes[1170]);
    tranif1 (nodes[1073], nodes[1326],  nodes[943]);
    tranif1 (nodes[7], nodes[558],  nodes[466]);
    tranif1 (nodes[471], nodes[657],  nodes[466]);
    tranif1 (nodes[558], nodes[384],  nodes[1258]);
    tranif1 (nodes[558], nodes[22],  nodes[193]);
    tranif1 (nodes[558], nodes[997],  nodes[289]);
    tranif1 (nodes[521], nodes[1358],  nodes[943]);
    tranif1 (nodes[1444], nodes[558],  nodes[318]);
    tranif1 (nodes[657], nodes[1443],  nodes[1545]);
    tranif1 (nodes[428], nodes[644],  nodes[710]);
    tranif1 (nodes[519], nodes[558],  nodes[1171]);
    tranif1 (nodes[558], nodes[1089],  nodes[1574]);
    tranif1 (nodes[1219], nodes[558],  nodes[776]);
    tranif1 (nodes[558], nodes[184],  nodes[305]);
    tranif1 (nodes[558], nodes[1079],  nodes[1411]);
    tranif1 (nodes[247], nodes[558],  nodes[849]);
    tranif1 (nodes[558], nodes[1211],  nodes[862]);
    tranif1 (nodes[1024], nodes[558],  nodes[94]);
    tranif1 (nodes[877], nodes[558],  nodes[933]);
    tranif1 (nodes[1406], nodes[1657],  nodes[523]);
    tranif1 (nodes[1659], nodes[875],  nodes[523]);
    tranif1 (nodes[743], nodes[558],  nodes[523]);
    tranif1 (nodes[513], nodes[558],  nodes[1646]);
    tranif1 (nodes[558], nodes[708],  nodes[1230]);
    tranif1 (nodes[549], nodes[657],  nodes[1230]);
    tranif1 (nodes[1398], nodes[304],  nodes[59]);
    tranif1 (nodes[957], nodes[143],  nodes[59]);
    tranif1 (nodes[1654], nodes[558],  nodes[947]);
    tranif1 (nodes[232], nodes[558],  nodes[377]);
    tranif1 (nodes[332], nodes[413],  nodes[1468]);
    tranif1 (nodes[558], nodes[1622],  nodes[758]);
    tranif1 (nodes[1190], nodes[558],  nodes[81]);
    tranif1 (nodes[1182], nodes[1300],  nodes[943]);
    tranif1 (nodes[1544], nodes[922],  nodes[270]);
    tranif1 (nodes[558], nodes[1115],  nodes[270]);
    tranif1 (nodes[110], nodes[558],  nodes[1691]);
    tranif1 (nodes[1023], nodes[558],  nodes[1691]);
    tranif1 (nodes[558], nodes[723],  nodes[868]);
    tranif1 (nodes[558], nodes[794],  nodes[746]);
    tranif1 (nodes[558], nodes[288],  nodes[746]);
    tranif1 (nodes[558], nodes[1681],  nodes[546]);
    tranif1 (nodes[558], nodes[1270],  nodes[43]);
    tranif1 (nodes[558], nodes[898],  nodes[1247]);
    tranif1 (nodes[1626], nodes[558],  nodes[119]);
    tranif1 (nodes[1197], nodes[1390],  nodes[500]);
    tranif1 (nodes[174], nodes[558],  nodes[500]);
    tranif1 (nodes[558], nodes[690],  nodes[188]);
    tranif1 (nodes[1040], nodes[782],  nodes[1303]);
    tranif1 (nodes[558], nodes[212],  nodes[1160]);
    tranif1 (nodes[819], nodes[558],  nodes[449]);
    tranif1 (nodes[558], nodes[457],  nodes[1302]);
    tranif1 (nodes[1015], nodes[558],  nodes[1033]);
    tranif1 (nodes[1299], nodes[1611],  nodes[414]);
    tranif1 (nodes[1188], nodes[305],  nodes[325]);
    tranif1 (nodes[55], nodes[11],  nodes[943]);
    tranif1 (nodes[1069], nodes[558],  nodes[1274]);
    tranif1 (nodes[1274], nodes[913],  nodes[710]);
    tranif1 (nodes[604], nodes[558],  nodes[1311]);
    tranif1 (nodes[298], nodes[558],  nodes[23]);
    tranif1 (nodes[1501], nodes[657],  nodes[23]);
    tranif1 (nodes[558], nodes[1093],  nodes[968]);
    tranif1 (nodes[1020], nodes[1705],  nodes[943]);
    tranif1 (nodes[781], nodes[558],  nodes[199]);
    tranif1 (nodes[1422], nodes[558],  nodes[199]);
    tranif1 (nodes[118], nodes[558],  nodes[334]);
    tranif1 (nodes[558], nodes[619],  nodes[700]);
    tranif1 (nodes[1090], nodes[558],  nodes[157]);
    tranif1 (nodes[1467], nodes[558],  nodes[1129]);
    tranif1 (nodes[736], nodes[657],  nodes[1633]);
    tranif1 (nodes[736], nodes[657],  nodes[1633]);
    tranif1 (nodes[736], nodes[657],  nodes[1633]);
    tranif1 (nodes[736], nodes[657],  nodes[1633]);
    tranif1 (nodes[736], nodes[657],  nodes[1633]);
    tranif1 (nodes[558], nodes[1556],  nodes[901]);
    tranif1 (nodes[558], nodes[867],  nodes[901]);
    tranif1 (nodes[558], nodes[1220],  nodes[647]);
    tranif1 (nodes[558], nodes[821],  nodes[1067]);
    tranif1 (nodes[1320], nodes[541],  nodes[943]);
    tranif1 (nodes[916], nodes[1409],  nodes[710]);
    tranif1 (nodes[862], nodes[558],  nodes[666]);
    tranif1 (nodes[558], nodes[283],  nodes[1323]);
    tranif1 (nodes[1206], nodes[558],  nodes[535]);
    tranif1 (nodes[558], nodes[1215],  nodes[1185]);
    tranif1 (nodes[558], nodes[1433],  nodes[201]);
    tranif1 (nodes[558], nodes[1200],  nodes[493]);
    tranif1 (nodes[744], nodes[558],  nodes[493]);
    tranif1 (nodes[967], nodes[558],  nodes[636]);
    tranif1 (nodes[657], nodes[268],  nodes[855]);
    tranif1 (nodes[657], nodes[268],  nodes[855]);
    tranif1 (nodes[657], nodes[268],  nodes[855]);
    tranif1 (nodes[657], nodes[268],  nodes[855]);
    tranif1 (nodes[657], nodes[268],  nodes[855]);
    tranif1 (nodes[1343], nodes[558],  nodes[248]);
    tranif1 (nodes[558], nodes[202],  nodes[646]);
    tranif1 (nodes[881], nodes[558],  nodes[943]);
    tranif1 (nodes[739], nodes[1080],  nodes[1056]);
    tranif1 (nodes[657], nodes[1539],  nodes[943]);
    tranif1 (nodes[558], nodes[631],  nodes[878]);
    tranif1 (nodes[1185], nodes[558],  nodes[916]);
    tranif1 (nodes[272], nodes[558],  nodes[967]);
    tranif1 (nodes[1333], nodes[80],  nodes[943]);
    tranif1 (nodes[558], nodes[571],  nodes[1671]);
    tranif1 (nodes[302], nodes[558],  nodes[1671]);
    tranif1 (nodes[558], nodes[1019],  nodes[1671]);
    tranif1 (nodes[1294], nodes[558],  nodes[1671]);
    tranif1 (nodes[558], nodes[1306],  nodes[1516]);
    tranif1 (nodes[1306], nodes[558],  nodes[1516]);
    tranif1 (nodes[558], nodes[1306],  nodes[1516]);
    tranif1 (nodes[1468], nodes[558],  nodes[196]);
    tranif1 (nodes[1058], nodes[558],  nodes[271]);
    tranif1 (nodes[24], nodes[1039],  nodes[710]);
    tranif1 (nodes[1649], nodes[558],  nodes[857]);
    tranif1 (nodes[1377], nodes[558],  nodes[857]);
    tranif1 (nodes[190], nodes[1101],  nodes[943]);
    tranif1 (nodes[558], nodes[412],  nodes[164]);
    tranif1 (nodes[20], nodes[993],  nodes[943]);
    tranif1 (nodes[558], nodes[726],  nodes[0]);
    tranif1 (nodes[558], nodes[1412],  nodes[1455]);
    tranif1 (nodes[1296], nodes[558],  nodes[1346]);
    tranif1 (nodes[657], nodes[359],  nodes[1346]);
    tranif1 (nodes[1455], nodes[558],  nodes[1324]);
    tranif1 (nodes[1001], nodes[765],  nodes[214]);
    tranif1 (nodes[104], nodes[558],  nodes[847]);
    tranif1 (nodes[1455], nodes[558],  nodes[1243]);
    tranif1 (nodes[148], nodes[558],  nodes[676]);
    tranif1 (nodes[558], nodes[148],  nodes[676]);
    tranif1 (nodes[148], nodes[558],  nodes[676]);
    tranif1 (nodes[558], nodes[148],  nodes[676]);
    tranif1 (nodes[148], nodes[558],  nodes[676]);
    tranif1 (nodes[148], nodes[558],  nodes[676]);
    tranif1 (nodes[148], nodes[558],  nodes[676]);
    tranif1 (nodes[1241], nodes[558],  nodes[748]);
    tranif1 (nodes[657], nodes[399],  nodes[1296]);
    tranif1 (nodes[267], nodes[558],  nodes[785]);
    tranif1 (nodes[657], nodes[353],  nodes[1028]);
    tranif1 (nodes[450], nodes[558],  nodes[1159]);
    tranif1 (nodes[558], nodes[1578],  nodes[1431]);
    tranif1 (nodes[558], nodes[1215],  nodes[238]);
    tranif1 (nodes[558], nodes[801],  nodes[969]);
    tranif1 (nodes[585], nodes[558],  nodes[232]);
    tranif1 (nodes[558], nodes[1704],  nodes[232]);
    tranif1 (nodes[1316], nodes[558],  nodes[232]);
    tranif1 (nodes[1069], nodes[1177],  nodes[943]);
    tranif1 (nodes[558], nodes[1315],  nodes[1429]);
    tranif1 (nodes[558], nodes[381],  nodes[1429]);
    tranif1 (nodes[1045], nodes[1442],  nodes[943]);
    tranif1 (nodes[1134], nodes[558],  nodes[1481]);
    tranif1 (nodes[357], nodes[728],  nodes[943]);
    tranif1 (nodes[160], nodes[558],  nodes[781]);
    tranif1 (nodes[912], nodes[558],  nodes[1481]);
    tranif1 (nodes[385], nodes[1652],  nodes[943]);
    tranif1 (nodes[558], nodes[1005],  nodes[558]);
    tranif1 (nodes[558], nodes[470],  nodes[646]);
    tranif1 (nodes[99], nodes[1194],  nodes[943]);
    tranif1 (nodes[558], nodes[556],  nodes[727]);
    tranif1 (nodes[558], nodes[368],  nodes[932]);
    tranif1 (nodes[1352], nodes[558],  nodes[932]);
    tranif1 (nodes[558], nodes[291],  nodes[1121]);
    tranif1 (nodes[733], nodes[558],  nodes[981]);
    tranif1 (nodes[66], nodes[107],  nodes[943]);
    tranif1 (nodes[657], nodes[475],  nodes[1143]);
    tranif1 (nodes[1677], nodes[558],  nodes[1143]);
    tranif1 (nodes[999], nodes[558],  nodes[1143]);
    tranif1 (nodes[394], nodes[957],  nodes[943]);
    tranif1 (nodes[558], nodes[1506],  nodes[1285]);
    tranif1 (nodes[1122], nodes[1510],  nodes[1285]);
    tranif1 (nodes[1175], nodes[558],  nodes[1447]);
    tranif1 (nodes[558], nodes[808],  nodes[1327]);
    tranif1 (nodes[558], nodes[1154],  nodes[959]);
    tranif1 (nodes[1493], nodes[558],  nodes[171]);
    tranif1 (nodes[1493], nodes[558],  nodes[171]);
    tranif1 (nodes[1493], nodes[558],  nodes[171]);
    tranif1 (nodes[1493], nodes[558],  nodes[171]);
    tranif1 (nodes[1686], nodes[1475],  nodes[345]);
    tranif1 (nodes[1097], nodes[558],  nodes[345]);
    tranif1 (nodes[767], nodes[558],  nodes[1138]);
    tranif1 (nodes[240], nodes[1387],  nodes[710]);
    tranif1 (nodes[1193], nodes[558],  nodes[815]);
    tranif1 (nodes[1065], nodes[558],  nodes[1292]);
    tranif1 (nodes[558], nodes[667],  nodes[829]);
    tranif1 (nodes[558], nodes[1434],  nodes[98]);
    tranif1 (nodes[558], nodes[830],  nodes[1505]);
    tranif1 (nodes[558], nodes[1030],  nodes[757]);
    tranif1 (nodes[671], nodes[1718],  nodes[710]);
    tranif1 (nodes[558], nodes[1130],  nodes[192]);
    tranif1 (nodes[1069], nodes[558],  nodes[1024]);
    tranif1 (nodes[1176], nodes[1231],  nodes[943]);
    tranif1 (nodes[558], nodes[1429],  nodes[1062]);
    tranif1 (nodes[358], nodes[558],  nodes[1171]);
    tranif1 (nodes[1090], nodes[558],  nodes[1222]);
    tranif1 (nodes[1717], nodes[558],  nodes[382]);
    tranif1 (nodes[54], nodes[1216],  nodes[1186]);
    tranif1 (nodes[482], nodes[1459],  nodes[336]);
    tranif1 (nodes[558], nodes[159],  nodes[558]);
    tranif1 (nodes[221], nodes[558],  nodes[1579]);
    tranif1 (nodes[892], nodes[1119],  nodes[1042]);
    tranif1 (nodes[558], nodes[374],  nodes[1591]);
    tranif1 (nodes[1302], nodes[439],  nodes[1042]);
    tranif1 (nodes[833], nodes[77],  nodes[1042]);
    tranif1 (nodes[558], nodes[279],  nodes[507]);
    tranif1 (nodes[1082], nodes[186],  nodes[507]);
    tranif1 (nodes[1266], nodes[961],  nodes[710]);
    tranif1 (nodes[1486], nodes[558],  nodes[200]);
    tranif1 (nodes[1367], nodes[293],  nodes[200]);
    tranif1 (nodes[57], nodes[558],  nodes[200]);
    tranif1 (nodes[558], nodes[1501],  nodes[353]);
    tranif1 (nodes[558], nodes[1501],  nodes[353]);
    tranif1 (nodes[1509], nodes[952],  nodes[943]);
    tranif1 (nodes[558], nodes[97],  nodes[222]);
    tranif1 (nodes[558], nodes[1245],  nodes[938]);
    tranif1 (nodes[1644], nodes[558],  nodes[99]);
    tranif1 (nodes[558], nodes[1666],  nodes[108]);
    tranif1 (nodes[558], nodes[1446],  nodes[850]);
    tranif1 (nodes[558], nodes[430],  nodes[850]);
    tranif1 (nodes[1216], nodes[1169],  nodes[943]);
    tranif1 (nodes[529], nodes[588],  nodes[943]);
    tranif1 (nodes[657], nodes[483],  nodes[943]);
    tranif1 (nodes[657], nodes[121],  nodes[943]);
    tranif1 (nodes[14], nodes[558],  nodes[67]);
    tranif1 (nodes[297], nodes[558],  nodes[1032]);
    tranif1 (nodes[763], nodes[558],  nodes[1534]);
    tranif1 (nodes[657], nodes[1068],  nodes[1534]);
    tranif1 (nodes[558], nodes[1045],  nodes[69]);
    tranif1 (nodes[1322], nodes[1009],  nodes[36]);
    tranif1 (nodes[735], nodes[558],  nodes[36]);
    tranif1 (nodes[539], nodes[657],  nodes[417]);
    tranif1 (nodes[657], nodes[539],  nodes[417]);
    tranif1 (nodes[657], nodes[539],  nodes[417]);
    tranif1 (nodes[539], nodes[657],  nodes[417]);
    tranif1 (nodes[539], nodes[657],  nodes[417]);
    tranif1 (nodes[539], nodes[657],  nodes[417]);
    tranif1 (nodes[657], nodes[539],  nodes[417]);
    tranif1 (nodes[558], nodes[1211],  nodes[967]);
    tranif1 (nodes[558], nodes[1211],  nodes[967]);
    tranif1 (nodes[558], nodes[1211],  nodes[1286]);
    tranif1 (nodes[1612], nodes[558],  nodes[690]);
    tranif1 (nodes[804], nodes[558],  nodes[690]);
    tranif1 (nodes[558], nodes[1311],  nodes[690]);
    tranif1 (nodes[558], nodes[492],  nodes[690]);
    tranif1 (nodes[558], nodes[1259],  nodes[690]);
    tranif1 (nodes[354], nodes[558],  nodes[690]);
    tranif1 (nodes[341], nodes[558],  nodes[690]);
    tranif1 (nodes[461], nodes[558],  nodes[690]);
    tranif1 (nodes[352], nodes[558],  nodes[690]);
    tranif1 (nodes[1589], nodes[558],  nodes[690]);
    tranif1 (nodes[558], nodes[1569],  nodes[690]);
    tranif1 (nodes[558], nodes[281],  nodes[690]);
    tranif1 (nodes[710], nodes[657],  nodes[1399]);
    tranif1 (nodes[558], nodes[321],  nodes[398]);
    tranif1 (nodes[558], nodes[692],  nodes[43]);
    tranif1 (nodes[558], nodes[620],  nodes[1293]);
    tranif1 (nodes[558], nodes[1122],  nodes[936]);
    tranif1 (nodes[558], nodes[1194],  nodes[348]);
    tranif1 (nodes[558], nodes[988],  nodes[350]);
    tranif1 (nodes[875], nodes[558],  nodes[743]);
    tranif1 (nodes[609], nodes[545],  nodes[743]);
    tranif1 (nodes[1547], nodes[558],  nodes[743]);
    tranif1 (nodes[1694], nodes[558],  nodes[890]);
    tranif1 (nodes[1001], nodes[1539],  nodes[140]);
    tranif1 (nodes[13], nodes[1336],  nodes[140]);
    tranif1 (nodes[54], nodes[64],  nodes[325]);
    tranif1 (nodes[54], nodes[407],  nodes[140]);
    tranif1 (nodes[558], nodes[38],  nodes[710]);
    tranif1 (nodes[1247], nodes[558],  nodes[710]);
    tranif1 (nodes[558], nodes[882],  nodes[1252]);
    tranif1 (nodes[1405], nodes[1160],  nodes[140]);
    tranif1 (nodes[1188], nodes[315],  nodes[140]);
    tranif1 (nodes[1287], nodes[1651],  nodes[140]);
    tranif1 (nodes[970], nodes[233],  nodes[761]);
    tranif1 (nodes[762], nodes[558],  nodes[761]);
    tranif1 (nodes[1372], nodes[558],  nodes[1201]);
    tranif1 (nodes[1293], nodes[558],  nodes[840]);
    tranif1 (nodes[558], nodes[1439],  nodes[115]);
    tranif1 (nodes[1072], nodes[558],  nodes[97]);
    tranif1 (nodes[769], nodes[558],  nodes[97]);
    tranif1 (nodes[1170], nodes[558],  nodes[755]);
    tranif1 (nodes[102], nodes[657],  nodes[834]);
    tranif1 (nodes[558], nodes[129],  nodes[75]);
    tranif1 (nodes[558], nodes[1571],  nodes[142]);
    tranif1 (nodes[165], nodes[427],  nodes[142]);
    tranif1 (nodes[957], nodes[1628],  nodes[574]);
    tranif1 (nodes[250], nodes[841],  nodes[574]);
    tranif1 (nodes[740], nodes[681],  nodes[574]);
    tranif1 (nodes[1071], nodes[350],  nodes[574]);
    tranif1 (nodes[296], nodes[1063],  nodes[574]);
    tranif1 (nodes[477], nodes[277],  nodes[574]);
    tranif1 (nodes[722], nodes[336],  nodes[574]);
    tranif1 (nodes[1318], nodes[304],  nodes[574]);
    tranif1 (nodes[569], nodes[1205],  nodes[233]);
    tranif1 (nodes[657], nodes[1282],  nodes[943]);
    tranif1 (nodes[887], nodes[657],  nodes[1191]);
    tranif1 (nodes[887], nodes[657],  nodes[1191]);
    tranif1 (nodes[887], nodes[657],  nodes[1191]);
    tranif1 (nodes[887], nodes[657],  nodes[1191]);
    tranif1 (nodes[709], nodes[558],  nodes[1499]);
    tranif1 (nodes[1201], nodes[657],  nodes[1499]);
    tranif1 (nodes[558], nodes[929],  nodes[1549]);
    tranif1 (nodes[558], nodes[414],  nodes[943]);
    tranif1 (nodes[558], nodes[898],  nodes[943]);
    tranif1 (nodes[132], nodes[558],  nodes[31]);
    tranif1 (nodes[558], nodes[1583],  nodes[918]);
    tranif1 (nodes[112], nodes[558],  nodes[336]);
    tranif1 (nodes[558], nodes[1110],  nodes[756]);
    tranif1 (nodes[1108], nodes[146],  nodes[1331]);
    tranif1 (nodes[991], nodes[929],  nodes[1331]);
    tranif1 (nodes[1473], nodes[1618],  nodes[1331]);
    tranif1 (nodes[1302], nodes[1654],  nodes[1331]);
    tranif1 (nodes[1344], nodes[892],  nodes[1331]);
    tranif1 (nodes[1503], nodes[831],  nodes[1331]);
    tranif1 (nodes[833], nodes[326],  nodes[1331]);
    tranif1 (nodes[493], nodes[1592],  nodes[1331]);
    tranif1 (nodes[558], nodes[540],  nodes[369]);
    tranif1 (nodes[1685], nodes[1542],  nodes[1345]);
    tranif1 (nodes[558], nodes[1568],  nodes[1345]);
    tranif1 (nodes[558], nodes[795],  nodes[1649]);
    tranif1 (nodes[1533], nodes[1180],  nodes[710]);
    tranif1 (nodes[983], nodes[558],  nodes[1403]);
    tranif1 (nodes[580], nodes[558],  nodes[1268]);
    tranif1 (nodes[1545], nodes[657],  nodes[287]);
    tranif1 (nodes[1034], nodes[558],  nodes[287]);
    tranif1 (nodes[994], nodes[558],  nodes[287]);
    tranif1 (nodes[347], nodes[558],  nodes[219]);
    tranif1 (nodes[52], nodes[1150],  nodes[140]);
    tranif1 (nodes[1332], nodes[558],  nodes[984]);
    tranif1 (nodes[582], nodes[558],  nodes[610]);
    tranif1 (nodes[1001], nodes[1251],  nodes[801]);
    tranif1 (nodes[558], nodes[937],  nodes[1139]);
    tranif1 (nodes[526], nodes[1500],  nodes[943]);
    tranif1 (nodes[1405], nodes[658],  nodes[801]);
    tranif1 (nodes[558], nodes[603],  nodes[47]);
    tranif1 (nodes[1336], nodes[518],  nodes[801]);
    tranif1 (nodes[166], nodes[733],  nodes[801]);
    tranif1 (nodes[558], nodes[499],  nodes[49]);
    tranif1 (nodes[824], nodes[558],  nodes[579]);
    tranif1 (nodes[445], nodes[558],  nodes[862]);
    tranif1 (nodes[1185], nodes[558],  nodes[729]);
    tranif1 (nodes[1519], nodes[738],  nodes[710]);
    tranif1 (nodes[734], nodes[558],  nodes[1540]);
    tranif1 (nodes[657], nodes[1503],  nodes[943]);
    tranif1 (nodes[629], nodes[558],  nodes[50]);
    tranif1 (nodes[151], nodes[440],  nodes[943]);
    tranif1 (nodes[558], nodes[1716],  nodes[660]);
    tranif1 (nodes[558], nodes[1708],  nodes[660]);
    tranif1 (nodes[256], nodes[558],  nodes[594]);
    tranif1 (nodes[208], nodes[558],  nodes[39]);
    tranif1 (nodes[1349], nodes[558],  nodes[558]);
    tranif1 (nodes[26], nodes[927],  nodes[943]);
    tranif1 (nodes[558], nodes[1335],  nodes[628]);
    tranif1 (nodes[1698], nodes[657],  nodes[628]);
    tranif1 (nodes[460], nodes[616],  nodes[943]);
    tranif1 (nodes[1233], nodes[558],  nodes[895]);
    tranif1 (nodes[76], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[1658],  nodes[895]);
    tranif1 (nodes[786], nodes[558],  nodes[895]);
    tranif1 (nodes[1664], nodes[558],  nodes[895]);
    tranif1 (nodes[1612], nodes[558],  nodes[895]);
    tranif1 (nodes[784], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[244],  nodes[895]);
    tranif1 (nodes[558], nodes[1623],  nodes[895]);
    tranif1 (nodes[764], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[1311],  nodes[895]);
    tranif1 (nodes[558], nodes[324],  nodes[895]);
    tranif1 (nodes[558], nodes[857],  nodes[895]);
    tranif1 (nodes[1337], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[1355],  nodes[895]);
    tranif1 (nodes[558], nodes[787],  nodes[895]);
    tranif1 (nodes[575], nodes[558],  nodes[895]);
    tranif1 (nodes[1381], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[822],  nodes[895]);
    tranif1 (nodes[558], nodes[131],  nodes[895]);
    tranif1 (nodes[1086], nodes[558],  nodes[895]);
    tranif1 (nodes[1074], nodes[558],  nodes[895]);
    tranif1 (nodes[1246], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[0],  nodes[895]);
    tranif1 (nodes[594], nodes[558],  nodes[895]);
    tranif1 (nodes[1052], nodes[558],  nodes[895]);
    tranif1 (nodes[1589], nodes[558],  nodes[895]);
    tranif1 (nodes[446], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[309],  nodes[895]);
    tranif1 (nodes[558], nodes[53],  nodes[895]);
    tranif1 (nodes[558], nodes[1292],  nodes[895]);
    tranif1 (nodes[1155], nodes[558],  nodes[895]);
    tranif1 (nodes[1569], nodes[558],  nodes[895]);
    tranif1 (nodes[301], nodes[558],  nodes[895]);
    tranif1 (nodes[950], nodes[558],  nodes[895]);
    tranif1 (nodes[1710], nodes[558],  nodes[895]);
    tranif1 (nodes[558], nodes[1419],  nodes[895]);
    tranif1 (nodes[716], nodes[558],  nodes[681]);
    tranif1 (nodes[1503], nodes[72],  nodes[283]);
    tranif1 (nodes[558], nodes[693],  nodes[143]);
    tranif1 (nodes[558], nodes[1285],  nodes[143]);
    tranif1 (nodes[604], nodes[558],  nodes[1031]);
    tranif1 (nodes[1505], nodes[1455],  nodes[943]);
    tranif1 (nodes[558], nodes[1240],  nodes[1566]);
    tranif1 (nodes[863], nodes[657],  nodes[1566]);
    tranif1 (nodes[864], nodes[1507],  nodes[710]);
    tranif1 (nodes[558], nodes[996],  nodes[1133]);
    tranif1 (nodes[919], nodes[856],  nodes[1704]);
    tranif1 (nodes[558], nodes[835],  nodes[1704]);
    tranif1 (nodes[558], nodes[838],  nodes[581]);
    tranif1 (nodes[1563], nodes[11],  nodes[397]);
    tranif1 (nodes[558], nodes[134],  nodes[1557]);
    tranif1 (nodes[208], nodes[892],  nodes[283]);
    tranif1 (nodes[558], nodes[1130],  nodes[862]);
    tranif1 (nodes[315], nodes[657],  nodes[943]);
    tranif1 (nodes[558], nodes[133],  nodes[943]);
    tranif1 (nodes[558], nodes[161],  nodes[943]);
    tranif1 (nodes[332], nodes[558],  nodes[418]);
    tranif1 (nodes[276], nodes[740],  nodes[943]);
    tranif1 (nodes[1000], nodes[558],  nodes[1466]);
    tranif1 (nodes[558], nodes[753],  nodes[1257]);
    tranif1 (nodes[558], nodes[711],  nodes[1257]);
    tranif1 (nodes[569], nodes[558],  nodes[1257]);
    tranif1 (nodes[558], nodes[440],  nodes[24]);
    tranif1 (nodes[558], nodes[1025],  nodes[64]);
    tranif1 (nodes[1107], nodes[558],  nodes[58]);
    tranif1 (nodes[360], nodes[795],  nodes[943]);
    tranif1 (nodes[1554], nodes[679],  nodes[739]);
    tranif1 (nodes[479], nodes[558],  nodes[739]);
    tranif1 (nodes[1631], nodes[868],  nodes[943]);
    tranif1 (nodes[272], nodes[558],  nodes[0]);
    tranif1 (nodes[1349], nodes[657],  nodes[298]);
    tranif1 (nodes[1349], nodes[657],  nodes[298]);
    tranif1 (nodes[1349], nodes[657],  nodes[298]);
    tranif1 (nodes[1349], nodes[657],  nodes[298]);
    tranif1 (nodes[195], nodes[558],  nodes[659]);
    tranif1 (nodes[558], nodes[195],  nodes[659]);
    tranif1 (nodes[558], nodes[195],  nodes[659]);
    tranif1 (nodes[558], nodes[195],  nodes[659]);
    tranif1 (nodes[195], nodes[558],  nodes[659]);
    tranif1 (nodes[558], nodes[195],  nodes[659]);
    tranif1 (nodes[146], nodes[54],  nodes[1698]);
    tranif1 (nodes[929], nodes[1150],  nodes[1698]);
    tranif1 (nodes[1287], nodes[1618],  nodes[1698]);
    tranif1 (nodes[1654], nodes[1188],  nodes[1698]);
    tranif1 (nodes[1344], nodes[1405],  nodes[1698]);
    tranif1 (nodes[831], nodes[166],  nodes[1698]);
    tranif1 (nodes[1336], nodes[326],  nodes[1698]);
    tranif1 (nodes[1001], nodes[1592],  nodes[1698]);
    tranif1 (nodes[694], nodes[1282],  nodes[1468]);
    tranif1 (nodes[642], nodes[707],  nodes[943]);
    tranif1 (nodes[558], nodes[1722],  nodes[780]);
    tranif1 (nodes[1704], nodes[558],  nodes[379]);
    tranif1 (nodes[558], nodes[1512],  nodes[1125]);
    tranif1 (nodes[382], nodes[558],  nodes[1125]);
    tranif1 (nodes[558], nodes[1173],  nodes[1125]);
    tranif1 (nodes[558], nodes[1543],  nodes[1125]);
    tranif1 (nodes[558], nodes[76],  nodes[1125]);
    tranif1 (nodes[558], nodes[245],  nodes[1125]);
    tranif1 (nodes[558], nodes[786],  nodes[1125]);
    tranif1 (nodes[558], nodes[1664],  nodes[1125]);
    tranif1 (nodes[558], nodes[682],  nodes[1125]);
    tranif1 (nodes[558], nodes[1482],  nodes[1125]);
    tranif1 (nodes[558], nodes[552],  nodes[1125]);
    tranif1 (nodes[558], nodes[1487],  nodes[1125]);
    tranif1 (nodes[558], nodes[764],  nodes[1125]);
    tranif1 (nodes[558], nodes[1057],  nodes[1125]);
    tranif1 (nodes[558], nodes[58],  nodes[1125]);
    tranif1 (nodes[558], nodes[1520],  nodes[1125]);
    tranif1 (nodes[558], nodes[1381],  nodes[1125]);
    tranif1 (nodes[558], nodes[257],  nodes[1125]);
    tranif1 (nodes[558], nodes[1324],  nodes[1125]);
    tranif1 (nodes[558], nodes[179],  nodes[1125]);
    tranif1 (nodes[131], nodes[558],  nodes[1125]);
    tranif1 (nodes[558], nodes[4],  nodes[1125]);
    tranif1 (nodes[558], nodes[1396],  nodes[1125]);
    tranif1 (nodes[558], nodes[167],  nodes[1125]);
    tranif1 (nodes[558], nodes[354],  nodes[1125]);
    tranif1 (nodes[558], nodes[1086],  nodes[1125]);
    tranif1 (nodes[558], nodes[1074],  nodes[1125]);
    tranif1 (nodes[273], nodes[558],  nodes[1125]);
    tranif1 (nodes[558], nodes[594],  nodes[1125]);
    tranif1 (nodes[558], nodes[677],  nodes[1125]);
    tranif1 (nodes[558], nodes[447],  nodes[1125]);
    tranif1 (nodes[558], nodes[1052],  nodes[1125]);
    tranif1 (nodes[791], nodes[558],  nodes[1125]);
    tranif1 (nodes[558], nodes[750],  nodes[1125]);
    tranif1 (nodes[558], nodes[932],  nodes[1125]);
    tranif1 (nodes[558], nodes[1589],  nodes[1125]);
    tranif1 (nodes[558], nodes[309],  nodes[1125]);
    tranif1 (nodes[558], nodes[1430],  nodes[1125]);
    tranif1 (nodes[558], nodes[1292],  nodes[1125]);
    tranif1 (nodes[558], nodes[1114],  nodes[1125]);
    tranif1 (nodes[558], nodes[1226],  nodes[1125]);
    tranif1 (nodes[558], nodes[1006],  nodes[1125]);
    tranif1 (nodes[558], nodes[1164],  nodes[1125]);
    tranif1 (nodes[558], nodes[950],  nodes[1125]);
    tranif1 (nodes[558], nodes[281],  nodes[1125]);
    tranif1 (nodes[558], nodes[1665],  nodes[1125]);
    tranif1 (nodes[558], nodes[607],  nodes[1125]);
    tranif1 (nodes[558], nodes[1419],  nodes[1125]);
    tranif1 (nodes[558], nodes[1050],  nodes[1125]);
    tranif1 (nodes[558], nodes[59],  nodes[1255]);
    tranif1 (nodes[558], nodes[1546],  nodes[781]);
    tranif1 (nodes[1457], nodes[558],  nodes[781]);
    tranif1 (nodes[1369], nodes[558],  nodes[897]);
    tranif1 (nodes[558], nodes[1508],  nodes[46]);
    tranif1 (nodes[1559], nodes[558],  nodes[530]);
    tranif1 (nodes[1632], nodes[558],  nodes[530]);
    tranif1 (nodes[510], nodes[558],  nodes[434]);
    tranif1 (nodes[558], nodes[414],  nodes[1247]);
    tranif1 (nodes[558], nodes[152],  nodes[630]);
    tranif1 (nodes[1572], nodes[558],  nodes[701]);
    tranif1 (nodes[193], nodes[558],  nodes[701]);
    tranif1 (nodes[558], nodes[1352],  nodes[335]);
    tranif1 (nodes[1156], nodes[558],  nodes[1696]);
    tranif1 (nodes[558], nodes[1156],  nodes[1696]);
    tranif1 (nodes[558], nodes[1156],  nodes[1696]);
    tranif1 (nodes[1156], nodes[558],  nodes[1696]);
    tranif1 (nodes[558], nodes[1156],  nodes[1696]);
    tranif1 (nodes[558], nodes[407],  nodes[229]);
    tranif1 (nodes[558], nodes[506],  nodes[192]);
    tranif1 (nodes[558], nodes[925],  nodes[517]);
    tranif1 (nodes[558], nodes[139],  nodes[934]);
    tranif1 (nodes[1711], nodes[1064],  nodes[943]);
    tranif1 (nodes[1443], nodes[657],  nodes[1545]);
    tranif1 (nodes[1181], nodes[648],  nodes[754]);
    tranif1 (nodes[558], nodes[1595],  nodes[754]);
    tranif1 (nodes[52], nodes[292],  nodes[48]);
    tranif1 (nodes[1178], nodes[590],  nodes[710]);
    tranif1 (nodes[775], nodes[558],  nodes[1128]);
    tranif1 (nodes[407], nodes[1670],  nodes[48]);
    tranif1 (nodes[558], nodes[617],  nodes[713]);
    tranif1 (nodes[558], nodes[676],  nodes[713]);
    tranif1 (nodes[1192], nodes[751],  nodes[943]);
    tranif1 (nodes[1639], nodes[657],  nodes[489]);
    tranif1 (nodes[1153], nodes[558],  nodes[489]);
    tranif1 (nodes[558], nodes[659],  nodes[489]);
    tranif1 (nodes[100], nodes[558],  nodes[1018]);
    tranif1 (nodes[558], nodes[1469],  nodes[1220]);
    tranif1 (nodes[778], nodes[558],  nodes[231]);
    tranif1 (nodes[368], nodes[558],  nodes[1430]);
    tranif1 (nodes[558], nodes[911],  nodes[877]);
    tranif1 (nodes[558], nodes[911],  nodes[877]);
    tranif1 (nodes[847], nodes[558],  nodes[300]);
    tranif1 (nodes[602], nodes[558],  nodes[133]);
    tranif1 (nodes[1263], nodes[657],  nodes[133]);
    tranif1 (nodes[558], nodes[1201],  nodes[709]);
    tranif1 (nodes[558], nodes[987],  nodes[1216]);
    tranif1 (nodes[1293], nodes[558],  nodes[318]);
    tranif1 (nodes[1075], nodes[558],  nodes[1393]);
    tranif1 (nodes[1007], nodes[558],  nodes[1704]);
    tranif1 (nodes[558], nodes[176],  nodes[236]);
    tranif1 (nodes[652], nodes[1551],  nodes[741]);
    tranif1 (nodes[1206], nodes[205],  nodes[741]);
    tranif1 (nodes[27], nodes[948],  nodes[741]);
    tranif1 (nodes[1301], nodes[49],  nodes[741]);
    tranif1 (nodes[1496], nodes[502],  nodes[741]);
    tranif1 (nodes[141], nodes[584],  nodes[741]);
    tranif1 (nodes[1722], nodes[1670],  nodes[741]);
    tranif1 (nodes[209], nodes[292],  nodes[741]);
    tranif1 (nodes[1411], nodes[515],  nodes[943]);
    tranif1 (nodes[558], nodes[616],  nodes[665]);
    tranif1 (nodes[315], nodes[558],  nodes[203]);
    tranif1 (nodes[1651], nodes[558],  nodes[203]);
    tranif1 (nodes[483], nodes[558],  nodes[203]);
    tranif1 (nodes[1160], nodes[558],  nodes[203]);
    tranif1 (nodes[558], nodes[550],  nodes[1228]);
    tranif1 (nodes[1539], nodes[558],  nodes[203]);
    tranif1 (nodes[13], nodes[558],  nodes[203]);
    tranif1 (nodes[558], nodes[1230],  nodes[360]);
    tranif1 (nodes[558], nodes[1118],  nodes[204]);
    tranif1 (nodes[1058], nodes[632],  nodes[1289]);
    tranif1 (nodes[198], nodes[558],  nodes[197]);
    tranif1 (nodes[198], nodes[558],  nodes[197]);
    tranif1 (nodes[1092], nodes[558],  nodes[888]);
    tranif1 (nodes[74], nodes[1675],  nodes[879]);
    tranif1 (nodes[1378], nodes[1609],  nodes[879]);
    tranif1 (nodes[1082], nodes[1692],  nodes[270]);
    tranif1 (nodes[558], nodes[1668],  nodes[407]);
    tranif1 (nodes[824], nodes[558],  nodes[487]);
    tranif1 (nodes[583], nodes[1432],  nodes[1068]);
    tranif1 (nodes[1621], nodes[96],  nodes[1068]);
    tranif1 (nodes[558], nodes[1619],  nodes[182]);
    tranif1 (nodes[1486], nodes[126],  nodes[943]);
    tranif1 (nodes[558], nodes[152],  nodes[788]);
    tranif1 (nodes[1492], nodes[558],  nodes[974]);
    tranif1 (nodes[558], nodes[378],  nodes[1357]);
    tranif1 (nodes[558], nodes[732],  nodes[1161]);
    tranif1 (nodes[1621], nodes[558],  nodes[1302]);
    tranif1 (nodes[182], nodes[558],  nodes[646]);
    tranif1 (nodes[347], nodes[558],  nodes[607]);
    tranif1 (nodes[1298], nodes[1267],  nodes[710]);
    tranif1 (nodes[42], nodes[558],  nodes[1613]);
    tranif1 (nodes[643], nodes[657],  nodes[1613]);
    tranif1 (nodes[1682], nodes[558],  nodes[901]);
    tranif1 (nodes[1362], nodes[558],  nodes[901]);
    tranif1 (nodes[378], nodes[940],  nodes[943]);
    tranif1 (nodes[187], nodes[558],  nodes[248]);
    tranif1 (nodes[1718], nodes[558],  nodes[248]);
    tranif1 (nodes[837], nodes[558],  nodes[1623]);
    tranif1 (nodes[657], nodes[1163],  nodes[747]);
    tranif1 (nodes[1715], nodes[558],  nodes[358]);
    tranif1 (nodes[208], nodes[1437],  nodes[438]);
    tranif1 (nodes[1630], nodes[72],  nodes[438]);
    tranif1 (nodes[1458], nodes[121],  nodes[438]);
    tranif1 (nodes[1299], nodes[1647],  nodes[438]);
    tranif1 (nodes[488], nodes[413],  nodes[438]);
    tranif1 (nodes[1282], nodes[976],  nodes[438]);
    tranif1 (nodes[481], nodes[1242],  nodes[438]);
    tranif1 (nodes[684], nodes[723],  nodes[438]);
    tranif1 (nodes[558], nodes[975],  nodes[854]);
    tranif1 (nodes[1500], nodes[558],  nodes[1345]);
    tranif1 (nodes[289], nodes[635],  nodes[943]);
    tranif1 (nodes[133], nodes[558],  nodes[1404]);
    tranif1 (nodes[1242], nodes[558],  nodes[1193]);
    tranif1 (nodes[1416], nodes[558],  nodes[833]);
    tranif1 (nodes[558], nodes[930],  nodes[1276]);
    tranif1 (nodes[558], nodes[930],  nodes[1276]);
    tranif1 (nodes[83], nodes[558],  nodes[1400]);
    tranif1 (nodes[558], nodes[611],  nodes[1509]);
    tranif1 (nodes[1507], nodes[558],  nodes[684]);
    tranif1 (nodes[657], nodes[43],  nodes[839]);
    tranif1 (nodes[536], nodes[484],  nodes[943]);
    tranif1 (nodes[558], nodes[6],  nodes[43]);
    tranif1 (nodes[1206], nodes[1539],  nodes[1235]);
    tranif1 (nodes[652], nodes[13],  nodes[1235]);
    tranif1 (nodes[1301], nodes[483],  nodes[1235]);
    tranif1 (nodes[27], nodes[1160],  nodes[1235]);
    tranif1 (nodes[141], nodes[315],  nodes[1235]);
    tranif1 (nodes[1496], nodes[1651],  nodes[1235]);
    tranif1 (nodes[209], nodes[52],  nodes[1235]);
    tranif1 (nodes[1722], nodes[407],  nodes[1235]);
    tranif1 (nodes[779], nodes[605],  nodes[1440]);
    tranif1 (nodes[700], nodes[558],  nodes[1201]);
    tranif1 (nodes[381], nodes[1062],  nodes[943]);
    tranif1 (nodes[558], nodes[1129],  nodes[710]);
    tranif1 (nodes[1352], nodes[558],  nodes[1642]);
    tranif1 (nodes[657], nodes[211],  nodes[1041]);
    tranif1 (nodes[211], nodes[657],  nodes[1041]);
    tranif1 (nodes[211], nodes[657],  nodes[1041]);
    tranif1 (nodes[211], nodes[657],  nodes[1041]);
    tranif1 (nodes[657], nodes[211],  nodes[1041]);
    tranif1 (nodes[558], nodes[1254],  nodes[178]);
    tranif1 (nodes[558], nodes[1195],  nodes[178]);
    tranif1 (nodes[1191], nodes[657],  nodes[178]);
    tranif1 (nodes[558], nodes[300],  nodes[389]);
    tranif1 (nodes[491], nodes[558],  nodes[1541]);
    tranif1 (nodes[657], nodes[437],  nodes[1541]);
    tranif1 (nodes[431], nodes[558],  nodes[943]);
    tranif1 (nodes[195], nodes[657],  nodes[1639]);
    tranif1 (nodes[657], nodes[1237],  nodes[475]);
    tranif1 (nodes[1072], nodes[558],  nodes[353]);
    tranif1 (nodes[1072], nodes[558],  nodes[353]);
    tranif1 (nodes[558], nodes[1189],  nodes[1008]);
    tranif1 (nodes[1511], nodes[558],  nodes[1008]);
    tranif1 (nodes[814], nodes[344],  nodes[410]);
    tranif1 (nodes[558], nodes[557],  nodes[410]);
    tranif1 (nodes[375], nodes[558],  nodes[308]);
    tranif1 (nodes[65], nodes[558],  nodes[308]);
    tranif1 (nodes[678], nodes[706],  nodes[943]);
    tranif1 (nodes[533], nodes[558],  nodes[561]);
    tranif1 (nodes[474], nodes[558],  nodes[410]);
    tranif1 (nodes[1608], nodes[558],  nodes[1423]);
    tranif1 (nodes[657], nodes[869],  nodes[1423]);
    tranif1 (nodes[836], nodes[168],  nodes[710]);
    tranif1 (nodes[558], nodes[1392],  nodes[1297]);
    tranif1 (nodes[1024], nodes[1699],  nodes[943]);
    tranif1 (nodes[1232], nodes[558],  nodes[364]);
    tranif1 (nodes[18], nodes[468],  nodes[710]);
    tranif1 (nodes[296], nodes[404],  nodes[59]);
    tranif1 (nodes[558], nodes[1649],  nodes[389]);
    tranif1 (nodes[1464], nodes[558],  nodes[1487]);
    tranif1 (nodes[277], nodes[1632],  nodes[59]);
    tranif1 (nodes[378], nodes[558],  nodes[18]);
    tranif1 (nodes[379], nodes[1480],  nodes[1570]);
    tranif1 (nodes[657], nodes[833],  nodes[943]);
    tranif1 (nodes[905], nodes[1681],  nodes[440]);
    tranif1 (nodes[576], nodes[213],  nodes[943]);
    tranif1 (nodes[537], nodes[862],  nodes[943]);
    tranif1 (nodes[158], nodes[789],  nodes[710]);
    tranif1 (nodes[558], nodes[1685],  nodes[1166]);
    tranif1 (nodes[558], nodes[1568],  nodes[1166]);
    tranif1 (nodes[855], nodes[558],  nodes[1660]);
    tranif1 (nodes[657], nodes[1100],  nodes[1660]);
    tranif1 (nodes[1712], nodes[558],  nodes[1134]);
    tranif1 (nodes[558], nodes[1006],  nodes[1050]);
    tranif1 (nodes[1594], nodes[656],  nodes[779]);
    tranif1 (nodes[1032], nodes[558],  nodes[297]);
    tranif1 (nodes[1344], nodes[558],  nodes[556]);
    tranif1 (nodes[1196], nodes[558],  nodes[1689]);
    tranif1 (nodes[826], nodes[558],  nodes[1315]);
    tranif1 (nodes[558], nodes[1202],  nodes[1265]);
    tranif1 (nodes[558], nodes[1334],  nodes[1265]);
    tranif1 (nodes[615], nodes[733],  nodes[943]);
    tranif1 (nodes[195], nodes[657],  nodes[1639]);
    tranif1 (nodes[558], nodes[63],  nodes[158]);
    tranif1 (nodes[1703], nodes[558],  nodes[1373]);
    tranif1 (nodes[395], nodes[558],  nodes[1373]);
    tranif1 (nodes[1639], nodes[558],  nodes[1153]);
    tranif1 (nodes[657], nodes[659],  nodes[1153]);
    tranif1 (nodes[558], nodes[761],  nodes[314]);
    tranif1 (nodes[1550], nodes[558],  nodes[781]);
    tranif1 (nodes[1269], nodes[967],  nodes[943]);
    tranif1 (nodes[1390], nodes[558],  nodes[1459]);
    tranif1 (nodes[174], nodes[558],  nodes[1459]);
    tranif1 (nodes[11], nodes[558],  nodes[1396]);
    tranif1 (nodes[327], nodes[199],  nodes[943]);
    tranif1 (nodes[338], nodes[252],  nodes[943]);
    tranif1 (nodes[1579], nodes[187],  nodes[710]);
    tranif1 (nodes[566], nodes[627],  nodes[710]);
    tranif1 (nodes[558], nodes[1186],  nodes[1247]);
    tranif1 (nodes[581], nodes[306],  nodes[943]);
    tranif1 (nodes[558], nodes[1564],  nodes[1157]);
    tranif1 (nodes[1374], nodes[558],  nodes[562]);
    tranif1 (nodes[558], nodes[1453],  nodes[1266]);
    tranif1 (nodes[657], nodes[195],  nodes[1639]);
    tranif1 (nodes[558], nodes[744],  nodes[1473]);
    tranif1 (nodes[314], nodes[558],  nodes[893]);
    tranif1 (nodes[1573], nodes[558],  nodes[1473]);
    tranif1 (nodes[558], nodes[662],  nodes[625]);
    tranif1 (nodes[1186], nodes[657],  nodes[625]);
    tranif1 (nodes[1172], nodes[558],  nodes[646]);
    tranif1 (nodes[464], nodes[558],  nodes[1284]);
    tranif1 (nodes[464], nodes[558],  nodes[1284]);
    tranif1 (nodes[464], nodes[558],  nodes[1284]);
    tranif1 (nodes[505], nodes[558],  nodes[1122]);
    tranif1 (nodes[433], nodes[558],  nodes[1122]);
    tranif1 (nodes[1213], nodes[558],  nodes[609]);
    tranif1 (nodes[657], nodes[1325],  nodes[97]);
    tranif1 (nodes[385], nodes[558],  nodes[604]);
    tranif1 (nodes[558], nodes[522],  nodes[1145]);
    tranif1 (nodes[5], nodes[558],  nodes[737]);
    tranif1 (nodes[1717], nodes[558],  nodes[1512]);
    tranif1 (nodes[17], nodes[554],  nodes[943]);
    tranif1 (nodes[1615], nodes[558],  nodes[940]);
    tranif1 (nodes[558], nodes[399],  nodes[359]);
    tranif1 (nodes[558], nodes[399],  nodes[359]);
    tranif1 (nodes[399], nodes[558],  nodes[359]);
    tranif1 (nodes[558], nodes[399],  nodes[359]);
    tranif1 (nodes[399], nodes[558],  nodes[359]);
    tranif1 (nodes[558], nodes[399],  nodes[359]);
    tranif1 (nodes[558], nodes[399],  nodes[359]);
    tranif1 (nodes[558], nodes[191],  nodes[790]);
    tranif1 (nodes[558], nodes[1107],  nodes[1204]);
    tranif1 (nodes[1638], nodes[558],  nodes[1591]);
    tranif1 (nodes[836], nodes[768],  nodes[821]);
    tranif1 (nodes[465], nodes[558],  nodes[206]);
    tranif1 (nodes[368], nodes[558],  nodes[528]);
    tranif1 (nodes[558], nodes[316],  nodes[1167]);
    tranif1 (nodes[143], nodes[558],  nodes[1167]);
    tranif1 (nodes[558], nodes[696],  nodes[217]);
    tranif1 (nodes[558], nodes[210],  nodes[234]);
    tranif1 (nodes[558], nodes[172],  nodes[234]);
    tranif1 (nodes[657], nodes[1633],  nodes[234]);
    tranif1 (nodes[558], nodes[1618],  nodes[419]);
    tranif1 (nodes[558], nodes[43],  nodes[710]);
    tranif1 (nodes[1247], nodes[558],  nodes[710]);
    tranif1 (nodes[558], nodes[1247],  nodes[710]);
    tranif1 (nodes[947], nodes[558],  nodes[162]);
    tranif1 (nodes[243], nodes[558],  nodes[991]);
    tranif1 (nodes[493], nodes[1535],  nodes[859]);
    tranif1 (nodes[833], nodes[235],  nodes[859]);
    tranif1 (nodes[558], nodes[60],  nodes[1576]);
    tranif1 (nodes[558], nodes[84],  nodes[1576]);
    tranif1 (nodes[558], nodes[271],  nodes[1576]);
    tranif1 (nodes[558], nodes[370],  nodes[1576]);
    tranif1 (nodes[558], nodes[1612],  nodes[1576]);
    tranif1 (nodes[558], nodes[784],  nodes[1576]);
    tranif1 (nodes[558], nodes[204],  nodes[1576]);
    tranif1 (nodes[558], nodes[804],  nodes[1576]);
    tranif1 (nodes[558], nodes[1311],  nodes[1576]);
    tranif1 (nodes[558], nodes[1428],  nodes[1576]);
    tranif1 (nodes[558], nodes[492],  nodes[1576]);
    tranif1 (nodes[558], nodes[1204],  nodes[1576]);
    tranif1 (nodes[558], nodes[1259],  nodes[1576]);
    tranif1 (nodes[558], nodes[342],  nodes[1576]);
    tranif1 (nodes[558], nodes[857],  nodes[1576]);
    tranif1 (nodes[558], nodes[712],  nodes[1576]);
    tranif1 (nodes[558], nodes[776],  nodes[1576]);
    tranif1 (nodes[558], nodes[1168],  nodes[1576]);
    tranif1 (nodes[558], nodes[1721],  nodes[1576]);
    tranif1 (nodes[558], nodes[487],  nodes[1576]);
    tranif1 (nodes[558], nodes[579],  nodes[1576]);
    tranif1 (nodes[558], nodes[1239],  nodes[1576]);
    tranif1 (nodes[558], nodes[285],  nodes[1576]);
    tranif1 (nodes[558], nodes[1524],  nodes[1576]);
    tranif1 (nodes[558], nodes[0],  nodes[1576]);
    tranif1 (nodes[558], nodes[1478],  nodes[1576]);
    tranif1 (nodes[558], nodes[1210],  nodes[1576]);
    tranif1 (nodes[558], nodes[461],  nodes[1576]);
    tranif1 (nodes[558], nodes[660],  nodes[1576]);
    tranif1 (nodes[558], nodes[1557],  nodes[1576]);
    tranif1 (nodes[558], nodes[259],  nodes[1576]);
    tranif1 (nodes[558], nodes[352],  nodes[1576]);
    tranif1 (nodes[558], nodes[446],  nodes[1576]);
    tranif1 (nodes[558], nodes[528],  nodes[1576]);
    tranif1 (nodes[558], nodes[904],  nodes[1576]);
    tranif1 (nodes[558], nodes[1569],  nodes[1576]);
    tranif1 (nodes[558], nodes[1710],  nodes[1576]);
    tranif1 (nodes[558], nodes[219],  nodes[1576]);
    tranif1 (nodes[558], nodes[1385],  nodes[1576]);
    tranif1 (nodes[391], nodes[1147],  nodes[710]);
    tranif1 (nodes[991], nodes[1432],  nodes[859]);
    tranif1 (nodes[1302], nodes[96],  nodes[859]);
    tranif1 (nodes[704], nodes[1473],  nodes[859]);
    tranif1 (nodes[1503], nodes[1678],  nodes[859]);
    tranif1 (nodes[892], nodes[1645],  nodes[859]);
    tranif1 (nodes[558], nodes[806],  nodes[558]);
    tranif1 (nodes[578], nodes[589],  nodes[943]);
    tranif1 (nodes[558], nodes[1586],  nodes[682]);
    tranif1 (nodes[994], nodes[768],  nodes[943]);
    tranif1 (nodes[426], nodes[1386],  nodes[1316]);
    tranif1 (nodes[558], nodes[914],  nodes[1316]);
    tranif1 (nodes[413], nodes[657],  nodes[943]);
    tranif1 (nodes[780], nodes[1229],  nodes[943]);
    tranif1 (nodes[558], nodes[41],  nodes[1441]);
    tranif1 (nodes[1695], nodes[1318],  nodes[1535]);
    tranif1 (nodes[1398], nodes[558],  nodes[1535]);
    tranif1 (nodes[20], nodes[558],  nodes[1316]);
    tranif1 (nodes[387], nodes[558],  nodes[853]);
    tranif1 (nodes[558], nodes[670],  nodes[519]);
    tranif1 (nodes[670], nodes[558],  nodes[519]);
    tranif1 (nodes[1302], nodes[723],  nodes[283]);
    tranif1 (nodes[991], nodes[976],  nodes[283]);
    tranif1 (nodes[1647], nodes[493],  nodes[283]);
    tranif1 (nodes[1481], nodes[558],  nodes[698]);
    tranif1 (nodes[558], nodes[1371],  nodes[846]);
    tranif1 (nodes[558], nodes[333],  nodes[1201]);
    tranif1 (nodes[558], nodes[228],  nodes[21]);
    tranif1 (nodes[48], nodes[657],  nodes[21]);
    tranif1 (nodes[1110], nodes[1530],  nodes[943]);
    tranif1 (nodes[558], nodes[765],  nodes[1123]);
    tranif1 (nodes[558], nodes[661],  nodes[1607]);
    tranif1 (nodes[558], nodes[1178],  nodes[1652]);
    tranif1 (nodes[1225], nodes[1121],  nodes[943]);
    tranif1 (nodes[558], nodes[549],  nodes[1247]);
    tranif1 (nodes[558], nodes[783],  nodes[655]);
    tranif1 (nodes[558], nodes[227],  nodes[540]);
    tranif1 (nodes[558], nodes[1263],  nodes[602]);
    tranif1 (nodes[464], nodes[1661],  nodes[710]);
    tranif1 (nodes[558], nodes[255],  nodes[611]);
    tranif1 (nodes[657], nodes[741],  nodes[611]);
    tranif1 (nodes[558], nodes[917],  nodes[248]);
    tranif1 (nodes[513], nodes[558],  nodes[954]);
    tranif1 (nodes[322], nodes[558],  nodes[1026]);
    tranif1 (nodes[657], nodes[171],  nodes[1026]);
    tranif1 (nodes[1082], nodes[455],  nodes[1051]);
    tranif1 (nodes[1249], nodes[626],  nodes[1200]);
    tranif1 (nodes[191], nodes[456],  nodes[943]);
    tranif1 (nodes[1455], nodes[558],  nodes[822]);
    tranif1 (nodes[558], nodes[918],  nodes[404]);
    tranif1 (nodes[558], nodes[142],  nodes[404]);
    tranif1 (nodes[1331], nodes[558],  nodes[943]);
    tranif1 (nodes[1698], nodes[558],  nodes[943]);
    tranif1 (nodes[1479], nodes[558],  nodes[842]);
    tranif1 (nodes[66], nodes[657],  nodes[842]);
    tranif1 (nodes[1140], nodes[657],  nodes[713]);
    tranif1 (nodes[558], nodes[1231],  nodes[1409]);
    tranif1 (nodes[558], nodes[11],  nodes[1228]);
    tranif1 (nodes[558], nodes[1135],  nodes[166]);
    tranif1 (nodes[558], nodes[1695],  nodes[1522]);
    tranif1 (nodes[1398], nodes[558],  nodes[1522]);
    tranif1 (nodes[86], nodes[364],  nodes[943]);
    tranif1 (nodes[558], nodes[1117],  nodes[70]);
    tranif1 (nodes[558], nodes[10],  nodes[1211]);
    tranif1 (nodes[1308], nodes[558],  nodes[637]);
    tranif1 (nodes[657], nodes[349],  nodes[1608]);
    tranif1 (nodes[431], nodes[807],  nodes[1599]);
    tranif1 (nodes[1698], nodes[558],  nodes[1335]);
    tranif1 (nodes[558], nodes[252],  nodes[1665]);
    tranif1 (nodes[1263], nodes[558],  nodes[1247]);
    tranif1 (nodes[1489], nodes[1308],  nodes[1314]);
    tranif1 (nodes[558], nodes[637],  nodes[1314]);
    tranif1 (nodes[819], nodes[558],  nodes[596]);
    tranif1 (nodes[658], nodes[558],  nodes[565]);
    tranif1 (nodes[1383], nodes[1678],  nodes[1068]);
    tranif1 (nodes[351], nodes[235],  nodes[1068]);
    tranif1 (nodes[423], nodes[1535],  nodes[1068]);
    tranif1 (nodes[558], nodes[1294],  nodes[1605]);
    tranif1 (nodes[558], nodes[1112],  nodes[927]);
    tranif1 (nodes[558], nodes[1449],  nodes[958]);
    tranif1 (nodes[777], nodes[871],  nodes[943]);
    tranif1 (nodes[835], nodes[1229],  nodes[919]);
    tranif1 (nodes[1538], nodes[1486],  nodes[919]);
    tranif1 (nodes[200], nodes[558],  nodes[919]);
    tranif1 (nodes[558], nodes[1655],  nodes[1211]);
    tranif1 (nodes[809], nodes[558],  nodes[1077]);
    tranif1 (nodes[1410], nodes[558],  nodes[1077]);
    tranif1 (nodes[1668], nodes[705],  nodes[710]);
    tranif1 (nodes[558], nodes[1211],  nodes[273]);
    tranif1 (nodes[1445], nodes[558],  nodes[1492]);
    tranif1 (nodes[1457], nodes[558],  nodes[1492]);
    tranif1 (nodes[525], nodes[558],  nodes[266]);
    tranif1 (nodes[188], nodes[558],  nodes[1357]);
    tranif1 (nodes[123], nodes[246],  nodes[710]);
    tranif1 (nodes[657], nodes[7],  nodes[1415]);
    tranif1 (nodes[413], nodes[558],  nodes[217]);
    tranif1 (nodes[813], nodes[558],  nodes[440]);
    tranif1 (nodes[1280], nodes[558],  nodes[335]);
    tranif1 (nodes[558], nodes[1549],  nodes[1234]);
    tranif1 (nodes[558], nodes[851],  nodes[302]);
    tranif1 (nodes[94], nodes[1650],  nodes[710]);
    tranif1 (nodes[506], nodes[1602],  nodes[943]);
    tranif1 (nodes[853], nodes[558],  nodes[770]);
    tranif1 (nodes[558], nodes[163],  nodes[249]);
    tranif1 (nodes[558], nodes[1704],  nodes[249]);
    tranif1 (nodes[558], nodes[890],  nodes[1]);
    tranif1 (nodes[1601], nodes[558],  nodes[1329]);
    tranif1 (nodes[382], nodes[558],  nodes[1329]);
    tranif1 (nodes[1173], nodes[558],  nodes[1329]);
    tranif1 (nodes[1233], nodes[558],  nodes[1329]);
    tranif1 (nodes[1543], nodes[558],  nodes[1329]);
    tranif1 (nodes[76], nodes[558],  nodes[1329]);
    tranif1 (nodes[1540], nodes[558],  nodes[1329]);
    tranif1 (nodes[558], nodes[245],  nodes[1329]);
    tranif1 (nodes[786], nodes[558],  nodes[1329]);
    tranif1 (nodes[1482], nodes[558],  nodes[1329]);
    tranif1 (nodes[370], nodes[558],  nodes[1329]);
    tranif1 (nodes[552], nodes[558],  nodes[1329]);
    tranif1 (nodes[784], nodes[558],  nodes[1329]);
    tranif1 (nodes[1623], nodes[558],  nodes[1329]);
    tranif1 (nodes[403], nodes[558],  nodes[1329]);
    tranif1 (nodes[558], nodes[1311],  nodes[1329]);
    tranif1 (nodes[1355], nodes[558],  nodes[1329]);
    tranif1 (nodes[257], nodes[558],  nodes[1329]);
    tranif1 (nodes[179], nodes[558],  nodes[1329]);
    tranif1 (nodes[1086], nodes[558],  nodes[1329]);
    tranif1 (nodes[487], nodes[558],  nodes[1329]);
    tranif1 (nodes[145], nodes[558],  nodes[1329]);
    tranif1 (nodes[1478], nodes[558],  nodes[1329]);
    tranif1 (nodes[558], nodes[1557],  nodes[1329]);
    tranif1 (nodes[517], nodes[558],  nodes[1329]);
    tranif1 (nodes[352], nodes[558],  nodes[1329]);
    tranif1 (nodes[750], nodes[558],  nodes[1329]);
    tranif1 (nodes[932], nodes[558],  nodes[1329]);
    tranif1 (nodes[309], nodes[558],  nodes[1329]);
    tranif1 (nodes[1569], nodes[558],  nodes[1329]);
    tranif1 (nodes[301], nodes[558],  nodes[1329]);
    tranif1 (nodes[941], nodes[558],  nodes[199]);
    tranif1 (nodes[558], nodes[25],  nodes[256]);
    tranif1 (nodes[1059], nodes[633],  nodes[943]);
    tranif1 (nodes[40], nodes[1575],  nodes[943]);
    tranif1 (nodes[558], nodes[1554],  nodes[61]);
    tranif1 (nodes[479], nodes[558],  nodes[61]);
    tranif1 (nodes[558], nodes[485],  nodes[85]);
    tranif1 (nodes[558], nodes[679],  nodes[479]);
    tranif1 (nodes[558], nodes[1088],  nodes[873]);
    tranif1 (nodes[134], nodes[558],  nodes[259]);
    tranif1 (nodes[558], nodes[444],  nodes[823]);
    tranif1 (nodes[558], nodes[1433],  nodes[840]);
    tranif1 (nodes[381], nodes[657],  nodes[1315]);
    tranif1 (nodes[523], nodes[949],  nodes[83]);
    tranif1 (nodes[1406], nodes[558],  nodes[83]);
    tranif1 (nodes[558], nodes[570],  nodes[1220]);
    tranif1 (nodes[264], nodes[799],  nodes[943]);
    tranif1 (nodes[264], nodes[1693],  nodes[943]);
    tranif1 (nodes[558], nodes[46],  nodes[992]);
    tranif1 (nodes[252], nodes[558],  nodes[301]);
    tranif1 (nodes[241], nodes[558],  nodes[745]);
    tranif1 (nodes[1446], nodes[558],  nodes[771]);
    tranif1 (nodes[465], nodes[430],  nodes[771]);
    tranif1 (nodes[766], nodes[474],  nodes[1184]);
    tranif1 (nodes[410], nodes[558],  nodes[1184]);
    tranif1 (nodes[558], nodes[1671],  nodes[1077]);
    tranif1 (nodes[1460], nodes[558],  nodes[1077]);
    tranif1 (nodes[558], nodes[811],  nodes[838]);
    tranif1 (nodes[26], nodes[558],  nodes[1112]);
    tranif1 (nodes[209], nodes[558],  nodes[113]);
    tranif1 (nodes[759], nodes[187],  nodes[710]);
    tranif1 (nodes[558], nodes[1687],  nodes[1108]);
    tranif1 (nodes[1035], nodes[558],  nodes[943]);
    tranif1 (nodes[1328], nodes[558],  nodes[541]);
    tranif1 (nodes[1150], nodes[872],  nodes[129]);
    tranif1 (nodes[558], nodes[587],  nodes[1283]);
    tranif1 (nodes[54], nodes[401],  nodes[129]);
    tranif1 (nodes[1109], nodes[558],  nodes[902]);
    tranif1 (nodes[1109], nodes[558],  nodes[902]);
    tranif1 (nodes[1289], nodes[558],  nodes[902]);
    tranif1 (nodes[558], nodes[1047],  nodes[830]);
    tranif1 (nodes[657], nodes[534],  nodes[830]);
    tranif1 (nodes[766], nodes[558],  nodes[1643]);
    tranif1 (nodes[558], nodes[1704],  nodes[1643]);
    tranif1 (nodes[410], nodes[558],  nodes[1643]);
    tranif1 (nodes[1587], nodes[558],  nodes[1077]);
    tranif1 (nodes[540], nodes[558],  nodes[1077]);
    tranif1 (nodes[1000], nodes[1408],  nodes[1044]);
    tranif1 (nodes[215], nodes[1379],  nodes[943]);
    tranif1 (nodes[345], nodes[1279],  nodes[986]);
    tranif1 (nodes[1108], nodes[1722],  nodes[247]);
    tranif1 (nodes[209], nodes[991],  nodes[247]);
    tranif1 (nodes[1496], nodes[1473],  nodes[247]);
    tranif1 (nodes[1302], nodes[141],  nodes[247]);
    tranif1 (nodes[892], nodes[27],  nodes[247]);
    tranif1 (nodes[1503], nodes[1301],  nodes[247]);
    tranif1 (nodes[652], nodes[833],  nodes[247]);
    tranif1 (nodes[1206], nodes[493],  nodes[247]);
    tranif1 (nodes[869], nodes[1128],  nodes[943]);
    tranif1 (nodes[558], nodes[772],  nodes[1674]);
    tranif1 (nodes[558], nodes[446],  nodes[909]);
    tranif1 (nodes[558], nodes[528],  nodes[909]);
    tranif1 (nodes[558], nodes[0],  nodes[909]);
    tranif1 (nodes[558], nodes[1210],  nodes[909]);
    tranif1 (nodes[558], nodes[1385],  nodes[909]);
    tranif1 (nodes[558], nodes[370],  nodes[909]);
    tranif1 (nodes[558], nodes[784],  nodes[909]);
    tranif1 (nodes[558], nodes[776],  nodes[909]);
    tranif1 (nodes[558], nodes[1168],  nodes[909]);
    tranif1 (nodes[1221], nodes[104],  nodes[943]);
    tranif1 (nodes[1186], nodes[558],  nodes[943]);
    tranif1 (nodes[558], nodes[1263],  nodes[943]);
    tranif1 (nodes[325], nodes[558],  nodes[943]);
    tranif1 (nodes[801], nodes[558],  nodes[943]);
    tranif1 (nodes[420], nodes[47],  nodes[710]);
    tranif1 (nodes[1706], nodes[558],  nodes[937]);
    tranif1 (nodes[1704], nodes[558],  nodes[937]);
    tranif1 (nodes[1345], nodes[558],  nodes[937]);
    tranif1 (nodes[558], nodes[717],  nodes[1132]);
    tranif1 (nodes[1380], nodes[666],  nodes[710]);
    tranif1 (nodes[558], nodes[334],  nodes[1382]);
    tranif1 (nodes[657], nodes[676],  nodes[617]);
    tranif1 (nodes[527], nodes[1474],  nodes[710]);
    tranif1 (nodes[558], nodes[1705],  nodes[630]);
    tranif1 (nodes[558], nodes[898],  nodes[1518]);
    tranif1 (nodes[558], nodes[1710],  nodes[996]);
    tranif1 (nodes[1601], nodes[558],  nodes[996]);
    tranif1 (nodes[382], nodes[558],  nodes[996]);
    tranif1 (nodes[1173], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[1233],  nodes[996]);
    tranif1 (nodes[558], nodes[1658],  nodes[996]);
    tranif1 (nodes[558], nodes[1664],  nodes[996]);
    tranif1 (nodes[558], nodes[1482],  nodes[996]);
    tranif1 (nodes[558], nodes[665],  nodes[996]);
    tranif1 (nodes[286], nodes[558],  nodes[996]);
    tranif1 (nodes[271], nodes[558],  nodes[996]);
    tranif1 (nodes[370], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[552],  nodes[996]);
    tranif1 (nodes[558], nodes[1612],  nodes[996]);
    tranif1 (nodes[558], nodes[1487],  nodes[996]);
    tranif1 (nodes[558], nodes[784],  nodes[996]);
    tranif1 (nodes[558], nodes[764],  nodes[996]);
    tranif1 (nodes[1582], nodes[558],  nodes[996]);
    tranif1 (nodes[1031], nodes[558],  nodes[996]);
    tranif1 (nodes[804], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[1311],  nodes[996]);
    tranif1 (nodes[558], nodes[1520],  nodes[996]);
    tranif1 (nodes[558], nodes[857],  nodes[996]);
    tranif1 (nodes[558], nodes[712],  nodes[996]);
    tranif1 (nodes[558], nodes[1337],  nodes[996]);
    tranif1 (nodes[1381], nodes[558],  nodes[996]);
    tranif1 (nodes[776], nodes[558],  nodes[996]);
    tranif1 (nodes[157], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[257],  nodes[996]);
    tranif1 (nodes[558], nodes[131],  nodes[996]);
    tranif1 (nodes[558], nodes[4],  nodes[996]);
    tranif1 (nodes[558], nodes[303],  nodes[996]);
    tranif1 (nodes[558], nodes[1721],  nodes[996]);
    tranif1 (nodes[1086], nodes[558],  nodes[996]);
    tranif1 (nodes[487], nodes[558],  nodes[996]);
    tranif1 (nodes[579], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[1239],  nodes[996]);
    tranif1 (nodes[558], nodes[0],  nodes[996]);
    tranif1 (nodes[558], nodes[1478],  nodes[996]);
    tranif1 (nodes[558], nodes[594],  nodes[996]);
    tranif1 (nodes[558], nodes[660],  nodes[996]);
    tranif1 (nodes[1557], nodes[558],  nodes[996]);
    tranif1 (nodes[259], nodes[558],  nodes[996]);
    tranif1 (nodes[1052], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[791],  nodes[996]);
    tranif1 (nodes[558], nodes[352],  nodes[996]);
    tranif1 (nodes[558], nodes[750],  nodes[996]);
    tranif1 (nodes[558], nodes[932],  nodes[996]);
    tranif1 (nodes[558], nodes[1589],  nodes[996]);
    tranif1 (nodes[446], nodes[558],  nodes[996]);
    tranif1 (nodes[528], nodes[558],  nodes[996]);
    tranif1 (nodes[309], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[1430],  nodes[996]);
    tranif1 (nodes[558], nodes[1292],  nodes[996]);
    tranif1 (nodes[558], nodes[1646],  nodes[996]);
    tranif1 (nodes[558], nodes[1114],  nodes[996]);
    tranif1 (nodes[558], nodes[1476],  nodes[996]);
    tranif1 (nodes[1226], nodes[558],  nodes[996]);
    tranif1 (nodes[1569], nodes[558],  nodes[996]);
    tranif1 (nodes[950], nodes[558],  nodes[996]);
    tranif1 (nodes[558], nodes[1050],  nodes[996]);
    tranif1 (nodes[558], nodes[1419],  nodes[996]);
    tranif1 (nodes[558], nodes[1164],  nodes[996]);
    tranif1 (nodes[558], nodes[995],  nodes[312]);
    tranif1 (nodes[742], nodes[854],  nodes[312]);
    tranif1 (nodes[558], nodes[1425],  nodes[988]);
    tranif1 (nodes[1382], nodes[1291],  nodes[710]);
    tranif1 (nodes[926], nodes[558],  nodes[717]);
    tranif1 (nodes[1087], nodes[558],  nodes[717]);
    tranif1 (nodes[1545], nodes[558],  nodes[1034]);
    tranif1 (nodes[657], nodes[994],  nodes[1034]);
    tranif1 (nodes[1410], nodes[558],  nodes[1690]);
    tranif1 (nodes[744], nodes[558],  nodes[1302]);
    tranif1 (nodes[558], nodes[1558],  nodes[40]);
    tranif1 (nodes[12], nodes[558],  nodes[40]);
    tranif1 (nodes[1016], nodes[558],  nodes[1282]);
    tranif1 (nodes[558], nodes[551],  nodes[393]);
    tranif1 (nodes[1085], nodes[596],  nodes[943]);
    tranif1 (nodes[685], nodes[1175],  nodes[943]);
    tranif1 (nodes[558], nodes[1312],  nodes[1291]);
    tranif1 (nodes[532], nodes[1013],  nodes[592]);
    tranif1 (nodes[1217], nodes[558],  nodes[592]);
    tranif1 (nodes[558], nodes[1510],  nodes[1021]);
    tranif1 (nodes[558], nodes[365],  nodes[809]);
    tranif1 (nodes[77], nodes[558],  nodes[90]);
    tranif1 (nodes[558], nodes[1454],  nodes[852]);
    tranif1 (nodes[558], nodes[260],  nodes[852]);
    tranif1 (nodes[1555], nodes[1107],  nodes[324]);
    tranif1 (nodes[1325], nodes[558],  nodes[769]);
    tranif1 (nodes[1072], nodes[657],  nodes[769]);
    tranif1 (nodes[1643], nodes[558],  nodes[900]);
    tranif1 (nodes[1393], nodes[1393],  nodes[147]);
    tranif1 (nodes[558], nodes[1393],  nodes[147]);
    tranif1 (nodes[558], nodes[1393],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[1393], nodes[558],  nodes[147]);
    tranif1 (nodes[558], nodes[1376],  nodes[1473]);
    tranif1 (nodes[125], nodes[558],  nodes[365]);
    tranif1 (nodes[558], nodes[363],  nodes[537]);
    tranif1 (nodes[558], nodes[731],  nodes[993]);
    tranif1 (nodes[1203], nodes[263],  nodes[753]);
    tranif1 (nodes[1629], nodes[558],  nodes[753]);
    tranif1 (nodes[558], nodes[827],  nodes[926]);
    tranif1 (nodes[339], nodes[632],  nodes[943]);
    tranif1 (nodes[108], nodes[558],  nodes[1364]);
    tranif1 (nodes[1666], nodes[657],  nodes[1364]);
    tranif1 (nodes[953], nodes[558],  nodes[425]);
    tranif1 (nodes[558], nodes[943],  nodes[1467]);
    tranif1 (nodes[558], nodes[943],  nodes[1467]);
    tranif1 (nodes[558], nodes[943],  nodes[1467]);
    tranif1 (nodes[943], nodes[558],  nodes[1467]);
    tranif1 (nodes[720], nodes[558],  nodes[56]);
    tranif1 (nodes[1494], nodes[558],  nodes[260]);
    tranif1 (nodes[558], nodes[1009],  nodes[735]);
    tranif1 (nodes[558], nodes[935],  nodes[1242]);
    tranif1 (nodes[146], nodes[558],  nodes[5]);
    tranif1 (nodes[558], nodes[438],  nodes[1462]);
    tranif1 (nodes[558], nodes[1544],  nodes[1115]);
    tranif1 (nodes[1658], nodes[558],  nodes[1394]);
    tranif1 (nodes[985], nodes[558],  nodes[1394]);
    tranif1 (nodes[1664], nodes[558],  nodes[1394]);
    tranif1 (nodes[682], nodes[558],  nodes[1394]);
    tranif1 (nodes[665], nodes[558],  nodes[1394]);
    tranif1 (nodes[286], nodes[558],  nodes[1394]);
    tranif1 (nodes[271], nodes[558],  nodes[1394]);
    tranif1 (nodes[1612], nodes[558],  nodes[1394]);
    tranif1 (nodes[1487], nodes[558],  nodes[1394]);
    tranif1 (nodes[244], nodes[558],  nodes[1394]);
    tranif1 (nodes[1520], nodes[558],  nodes[1394]);
    tranif1 (nodes[324], nodes[558],  nodes[1394]);
    tranif1 (nodes[712], nodes[558],  nodes[1394]);
    tranif1 (nodes[787], nodes[558],  nodes[1394]);
    tranif1 (nodes[575], nodes[558],  nodes[1394]);
    tranif1 (nodes[1466], nodes[558],  nodes[1394]);
    tranif1 (nodes[776], nodes[558],  nodes[1394]);
    tranif1 (nodes[822], nodes[558],  nodes[1394]);
    tranif1 (nodes[131], nodes[558],  nodes[1394]);
    tranif1 (nodes[1420], nodes[558],  nodes[1394]);
    tranif1 (nodes[4], nodes[558],  nodes[1394]);
    tranif1 (nodes[167], nodes[558],  nodes[1394]);
    tranif1 (nodes[303], nodes[558],  nodes[1394]);
    tranif1 (nodes[1504], nodes[558],  nodes[1394]);
    tranif1 (nodes[579], nodes[558],  nodes[1394]);
    tranif1 (nodes[0], nodes[558],  nodes[1394]);
    tranif1 (nodes[259], nodes[558],  nodes[1394]);
    tranif1 (nodes[528], nodes[558],  nodes[1394]);
    tranif1 (nodes[1430], nodes[558],  nodes[1394]);
    tranif1 (nodes[1646], nodes[558],  nodes[1394]);
    tranif1 (nodes[1155], nodes[558],  nodes[1394]);
    tranif1 (nodes[1476], nodes[558],  nodes[1394]);
    tranif1 (nodes[1226], nodes[558],  nodes[1394]);
    tranif1 (nodes[1164], nodes[558],  nodes[1394]);
    tranif1 (nodes[558], nodes[1497],  nodes[1438]);
    tranif1 (nodes[558], nodes[887],  nodes[1254]);
    tranif1 (nodes[887], nodes[558],  nodes[1254]);
    tranif1 (nodes[887], nodes[558],  nodes[1254]);
    tranif1 (nodes[887], nodes[558],  nodes[1254]);
    tranif1 (nodes[558], nodes[302],  nodes[540]);
    tranif1 (nodes[365], nodes[558],  nodes[540]);
    tranif1 (nodes[558], nodes[1294],  nodes[540]);
    tranif1 (nodes[506], nodes[558],  nodes[236]);
    tranif1 (nodes[558], nodes[1656],  nodes[1580]);
    tranif1 (nodes[558], nodes[1159],  nodes[1580]);
    tranif1 (nodes[1550], nodes[845],  nodes[1573]);
    tranif1 (nodes[558], nodes[959],  nodes[430]);
    tranif1 (nodes[166], nodes[578],  nodes[1263]);
    tranif1 (nodes[1336], nodes[1724],  nodes[1263]);
    tranif1 (nodes[574], nodes[558],  nodes[1256]);
    tranif1 (nodes[1287], nodes[1694],  nodes[1263]);
    tranif1 (nodes[1188], nodes[242],  nodes[1263]);
    tranif1 (nodes[1405], nodes[436],  nodes[1263]);
    tranif1 (nodes[520], nodes[558],  nodes[224]);
    tranif1 (nodes[37], nodes[657],  nodes[224]);
    tranif1 (nodes[831], nodes[558],  nodes[1719]);
    tranif1 (nodes[570], nodes[558],  nodes[1144]);
    tranif1 (nodes[558], nodes[1394],  nodes[1329]);
    tranif1 (nodes[879], nodes[558],  nodes[248]);
    tranif1 (nodes[538], nodes[558],  nodes[1599]);
    tranif1 (nodes[399], nodes[657],  nodes[1296]);
    tranif1 (nodes[1599], nodes[558],  nodes[103]);
    tranif1 (nodes[1577], nodes[1391],  nodes[943]);
    tranif1 (nodes[1255], nodes[558],  nodes[531]);
    tranif1 (nodes[59], nodes[657],  nodes[531]);
    tranif1 (nodes[298], nodes[657],  nodes[63]);
    tranif1 (nodes[999], nodes[668],  nodes[943]);
    tranif1 (nodes[907], nodes[1298],  nodes[821]);
    tranif1 (nodes[1404], nodes[1106],  nodes[943]);
    tranif1 (nodes[240], nodes[558],  nodes[498]);
    tranif1 (nodes[240], nodes[558],  nodes[498]);
    tranif1 (nodes[240], nodes[558],  nodes[498]);
    tranif1 (nodes[1464], nodes[558],  nodes[1612]);
    tranif1 (nodes[1649], nodes[558],  nodes[712]);
    tranif1 (nodes[1150], nodes[767],  nodes[801]);
    tranif1 (nodes[189], nodes[841],  nodes[1432]);
    tranif1 (nodes[155], nodes[558],  nodes[1432]);
    tranif1 (nodes[558], nodes[1186],  nodes[662]);
    tranif1 (nodes[33], nodes[558],  nodes[469]);
    tranif1 (nodes[558], nodes[86],  nodes[1232]);
    tranif1 (nodes[1676], nodes[558],  nodes[1232]);
    tranif1 (nodes[657], nodes[634],  nodes[1232]);
    tranif1 (nodes[1709], nodes[558],  nodes[1434]);
    tranif1 (nodes[1389], nodes[558],  nodes[752]);
    tranif1 (nodes[216], nodes[558],  nodes[681]);
    tranif1 (nodes[558], nodes[639],  nodes[130]);
    tranif1 (nodes[558], nodes[104],  nodes[275]);
    tranif1 (nodes[851], nodes[1515],  nodes[1019]);
    tranif1 (nodes[558], nodes[231],  nodes[1019]);
    tranif1 (nodes[558], nodes[1458],  nodes[731]);
    tranif1 (nodes[1120], nodes[558],  nodes[248]);
    tranif1 (nodes[2], nodes[1039],  nodes[248]);
    tranif1 (nodes[300], nodes[558],  nodes[342]);
    tranif1 (nodes[558], nodes[117],  nodes[1398]);
    tranif1 (nodes[1241], nodes[558],  nodes[1398]);
    tranif1 (nodes[1140], nodes[558],  nodes[617]);
    tranif1 (nodes[558], nodes[1295],  nodes[1527]);
    tranif1 (nodes[558], nodes[1515],  nodes[125]);
    tranif1 (nodes[90], nodes[558],  nodes[1625]);
    tranif1 (nodes[558], nodes[1379],  nodes[1476]);
    tranif1 (nodes[558], nodes[275],  nodes[1697]);
    tranif1 (nodes[595], nodes[558],  nodes[1168]);
    tranif1 (nodes[558], nodes[623],  nodes[143]);
    tranif1 (nodes[558], nodes[1347],  nodes[782]);
    tranif1 (nodes[558], nodes[934],  nodes[366]);
    tranif1 (nodes[72], nodes[622],  nodes[898]);
    tranif1 (nodes[208], nodes[900],  nodes[898]);
    tranif1 (nodes[1647], nodes[1611],  nodes[898]);
    tranif1 (nodes[1458], nodes[377],  nodes[898]);
    tranif1 (nodes[976], nodes[1022],  nodes[898]);
    tranif1 (nodes[488], nodes[1139],  nodes[898]);
    tranif1 (nodes[723], nodes[1359],  nodes[898]);
    tranif1 (nodes[481], nodes[655],  nodes[898]);
    tranif1 (nodes[166], nodes[483],  nodes[140]);
    tranif1 (nodes[121], nodes[618],  nodes[1468]);
    tranif1 (nodes[254], nodes[558],  nodes[483]);
    tranif1 (nodes[1038], nodes[558],  nodes[336]);
    tranif1 (nodes[1158], nodes[515],  nodes[1542]);
    tranif1 (nodes[1253], nodes[558],  nodes[1542]);
    tranif1 (nodes[558], nodes[984],  nodes[1247]);
    tranif1 (nodes[870], nodes[558],  nodes[576]);
    tranif1 (nodes[870], nodes[558],  nodes[576]);
    tranif1 (nodes[870], nodes[558],  nodes[576]);
    tranif1 (nodes[515], nodes[558],  nodes[1253]);
    tranif1 (nodes[160], nodes[558],  nodes[934]);
    tranif1 (nodes[558], nodes[1689],  nodes[837]);
    tranif1 (nodes[910], nodes[558],  nodes[590]);
    tranif1 (nodes[54], nodes[332],  nodes[1700]);
    tranif1 (nodes[423], nodes[558],  nodes[493]);
    tranif1 (nodes[774], nodes[974],  nodes[943]);
    tranif1 (nodes[968], nodes[934],  nodes[943]);
    tranif1 (nodes[415], nodes[1196],  nodes[943]);
    tranif1 (nodes[1688], nodes[680],  nodes[943]);
    tranif1 (nodes[558], nodes[106],  nodes[1528]);
    tranif1 (nodes[669], nodes[558],  nodes[303]);
    tranif1 (nodes[235], nodes[121],  nodes[437]);
    tranif1 (nodes[1535], nodes[1299],  nodes[437]);
    tranif1 (nodes[657], nodes[349],  nodes[1608]);
    tranif1 (nodes[1432], nodes[1282],  nodes[437]);
    tranif1 (nodes[1645], nodes[1437],  nodes[437]);
    tranif1 (nodes[1630], nodes[1678],  nodes[437]);
    tranif1 (nodes[1465], nodes[1126],  nodes[943]);
    tranif1 (nodes[96], nodes[684],  nodes[437]);
    tranif1 (nodes[899], nodes[19],  nodes[943]);
    tranif1 (nodes[1179], nodes[558],  nodes[725]);
    tranif1 (nodes[558], nodes[1286],  nodes[930]);
    tranif1 (nodes[718], nodes[558],  nodes[1005]);
    tranif1 (nodes[558], nodes[1591],  nodes[558]);
    tranif1 (nodes[978], nodes[1618],  nodes[943]);
    tranif1 (nodes[111], nodes[558],  nodes[945]);
    tranif1 (nodes[1123], nodes[304],  nodes[943]);
    tranif1 (nodes[558], nodes[896],  nodes[650]);
    tranif1 (nodes[558], nodes[1211],  nodes[1002]);
    tranif1 (nodes[299], nodes[1470],  nodes[1416]);
    tranif1 (nodes[558], nodes[152],  nodes[952]);
    tranif1 (nodes[272], nodes[558],  nodes[862]);
    tranif1 (nodes[1351], nodes[1717],  nodes[258]);
    tranif1 (nodes[1150], nodes[1709],  nodes[1263]);
    tranif1 (nodes[558], nodes[1228],  nodes[669]);
    tranif1 (nodes[558], nodes[1393],  nodes[558]);
    tranif1 (nodes[1252], nodes[1374],  nodes[943]);
    tranif1 (nodes[558], nodes[1483],  nodes[1627]);
    tranif1 (nodes[1084], nodes[558],  nodes[1627]);
    tranif1 (nodes[558], nodes[1707],  nodes[936]);
    tranif1 (nodes[558], nodes[388],  nodes[936]);
    tranif1 (nodes[1344], nodes[727],  nodes[943]);
    tranif1 (nodes[1265], nodes[558],  nodes[502]);
    tranif1 (nodes[1251], nodes[558],  nodes[1640]);
    tranif1 (nodes[420], nodes[558],  nodes[865]);
    tranif1 (nodes[558], nodes[645],  nodes[1032]);
    tranif1 (nodes[558], nodes[60],  nodes[1384]);
    tranif1 (nodes[558], nodes[1512],  nodes[1384]);
    tranif1 (nodes[558], nodes[382],  nodes[1384]);
    tranif1 (nodes[558], nodes[1173],  nodes[1384]);
    tranif1 (nodes[558], nodes[84],  nodes[1384]);
    tranif1 (nodes[558], nodes[1543],  nodes[1384]);
    tranif1 (nodes[558], nodes[76],  nodes[1384]);
    tranif1 (nodes[558], nodes[245],  nodes[1384]);
    tranif1 (nodes[558], nodes[786],  nodes[1384]);
    tranif1 (nodes[558], nodes[1664],  nodes[1384]);
    tranif1 (nodes[558], nodes[682],  nodes[1384]);
    tranif1 (nodes[558], nodes[1482],  nodes[1384]);
    tranif1 (nodes[558], nodes[271],  nodes[1384]);
    tranif1 (nodes[558], nodes[370],  nodes[1384]);
    tranif1 (nodes[558], nodes[552],  nodes[1384]);
    tranif1 (nodes[558], nodes[1612],  nodes[1384]);
    tranif1 (nodes[558], nodes[1487],  nodes[1384]);
    tranif1 (nodes[558], nodes[784],  nodes[1384]);
    tranif1 (nodes[558], nodes[1582],  nodes[1384]);
    tranif1 (nodes[558], nodes[804],  nodes[1384]);
    tranif1 (nodes[558], nodes[1311],  nodes[1384]);
    tranif1 (nodes[558], nodes[1428],  nodes[1384]);
    tranif1 (nodes[558], nodes[492],  nodes[1384]);
    tranif1 (nodes[558], nodes[1204],  nodes[1384]);
    tranif1 (nodes[558], nodes[1520],  nodes[1384]);
    tranif1 (nodes[558], nodes[1259],  nodes[1384]);
    tranif1 (nodes[558], nodes[342],  nodes[1384]);
    tranif1 (nodes[558], nodes[857],  nodes[1384]);
    tranif1 (nodes[558], nodes[712],  nodes[1384]);
    tranif1 (nodes[558], nodes[776],  nodes[1384]);
    tranif1 (nodes[558], nodes[157],  nodes[1384]);
    tranif1 (nodes[558], nodes[257],  nodes[1384]);
    tranif1 (nodes[558], nodes[1324],  nodes[1384]);
    tranif1 (nodes[558], nodes[179],  nodes[1384]);
    tranif1 (nodes[558], nodes[131],  nodes[1384]);
    tranif1 (nodes[558], nodes[4],  nodes[1384]);
    tranif1 (nodes[558], nodes[1396],  nodes[1384]);
    tranif1 (nodes[558], nodes[167],  nodes[1384]);
    tranif1 (nodes[558], nodes[1168],  nodes[1384]);
    tranif1 (nodes[558], nodes[1721],  nodes[1384]);
    tranif1 (nodes[558], nodes[1086],  nodes[1384]);
    tranif1 (nodes[558], nodes[1074],  nodes[1384]);
    tranif1 (nodes[558], nodes[487],  nodes[1384]);
    tranif1 (nodes[558], nodes[579],  nodes[1384]);
    tranif1 (nodes[558], nodes[1239],  nodes[1384]);
    tranif1 (nodes[558], nodes[1524],  nodes[1384]);
    tranif1 (nodes[558], nodes[0],  nodes[1384]);
    tranif1 (nodes[558], nodes[1478],  nodes[1384]);
    tranif1 (nodes[558], nodes[1210],  nodes[1384]);
    tranif1 (nodes[558], nodes[461],  nodes[1384]);
    tranif1 (nodes[558], nodes[660],  nodes[1384]);
    tranif1 (nodes[558], nodes[1557],  nodes[1384]);
    tranif1 (nodes[558], nodes[259],  nodes[1384]);
    tranif1 (nodes[558], nodes[791],  nodes[1384]);
    tranif1 (nodes[558], nodes[352],  nodes[1384]);
    tranif1 (nodes[558], nodes[750],  nodes[1384]);
    tranif1 (nodes[558], nodes[932],  nodes[1384]);
    tranif1 (nodes[558], nodes[446],  nodes[1384]);
    tranif1 (nodes[558], nodes[528],  nodes[1384]);
    tranif1 (nodes[558], nodes[1430],  nodes[1384]);
    tranif1 (nodes[558], nodes[1292],  nodes[1384]);
    tranif1 (nodes[558], nodes[1114],  nodes[1384]);
    tranif1 (nodes[558], nodes[1226],  nodes[1384]);
    tranif1 (nodes[558], nodes[1569],  nodes[1384]);
    tranif1 (nodes[558], nodes[1665],  nodes[1384]);
    tranif1 (nodes[558], nodes[1050],  nodes[1384]);
    tranif1 (nodes[558], nodes[1419],  nodes[1384]);
    tranif1 (nodes[558], nodes[1385],  nodes[1384]);
    tranif1 (nodes[558], nodes[1164],  nodes[1384]);
    tranif1 (nodes[558], nodes[1006],  nodes[1384]);
    tranif1 (nodes[45], nodes[1712],  nodes[943]);
    tranif1 (nodes[871], nodes[558],  nodes[1561]);
    tranif1 (nodes[558], nodes[726],  nodes[1210]);
    tranif1 (nodes[256], nodes[558],  nodes[1210]);
    tranif1 (nodes[1076], nodes[558],  nodes[1463]);
    tranif1 (nodes[147], nodes[657],  nodes[1463]);
    tranif1 (nodes[1711], nodes[558],  nodes[183]);
    tranif1 (nodes[1455], nodes[558],  nodes[257]);
    tranif1 (nodes[564], nodes[64],  nodes[943]);
    tranif1 (nodes[429], nodes[659],  nodes[943]);
    tranif1 (nodes[558], nodes[1209],  nodes[1213]);
    tranif1 (nodes[48], nodes[558],  nodes[228]);
    tranif1 (nodes[186], nodes[558],  nodes[1224]);
    tranif1 (nodes[1414], nodes[558],  nodes[495]);
    tranif1 (nodes[1441], nodes[558],  nodes[1277]);
    tranif1 (nodes[41], nodes[657],  nodes[1277]);
    tranif1 (nodes[781], nodes[558],  nodes[248]);
    tranif1 (nodes[781], nodes[558],  nodes[248]);
    tranif1 (nodes[558], nodes[930],  nodes[134]);
    tranif1 (nodes[558], nodes[467],  nodes[134]);
    tranif1 (nodes[67], nodes[449],  nodes[943]);
    tranif1 (nodes[558], nodes[1080],  nodes[811]);
    tranif1 (nodes[100], nodes[1205],  nodes[811]);
    tranif1 (nodes[657], nodes[991],  nodes[943]);
    tranif1 (nodes[1641], nodes[558],  nodes[809]);
    tranif1 (nodes[1547], nodes[1192],  nodes[609]);
    tranif1 (nodes[1264], nodes[1209],  nodes[609]);
    tranif1 (nodes[384], nodes[558],  nodes[1412]);
    tranif1 (nodes[558], nodes[62],  nodes[1349]);
    tranif1 (nodes[720], nodes[1338],  nodes[710]);
    tranif1 (nodes[1109], nodes[558],  nodes[1464]);
    tranif1 (nodes[703], nodes[227],  nodes[710]);
    tranif1 (nodes[657], nodes[166],  nodes[943]);
    tranif1 (nodes[181], nodes[548],  nodes[943]);
    tranif1 (nodes[1306], nodes[1095],  nodes[710]);
    tranif1 (nodes[43], nodes[558],  nodes[710]);
    tranif1 (nodes[839], nodes[558],  nodes[710]);
    tranif1 (nodes[507], nodes[558],  nodes[1049]);
    tranif1 (nodes[954], nodes[558],  nodes[338]);
    tranif1 (nodes[1522], nodes[1001],  nodes[549]);
    tranif1 (nodes[558], nodes[981],  nodes[615]);
    tranif1 (nodes[558], nodes[1260],  nodes[598]);
    tranif1 (nodes[328], nodes[558],  nodes[310]);
    tranif1 (nodes[558], nodes[494],  nodes[1539]);
    tranif1 (nodes[657], nodes[13],  nodes[943]);
    tranif1 (nodes[1299], nodes[657],  nodes[943]);
    tranif1 (nodes[558], nodes[501],  nodes[180]);
    tranif1 (nodes[558], nodes[976],  nodes[1102]);
    tranif1 (nodes[192], nodes[239],  nodes[1048]);
    tranif1 (nodes[1531], nodes[558],  nodes[184]);
    tranif1 (nodes[1485], nodes[1199],  nodes[943]);
    tranif1 (nodes[56], nodes[824],  nodes[943]);
    tranif1 (nodes[558], nodes[886],  nodes[943]);
    tranif1 (nodes[1307], nodes[524],  nodes[639]);
    tranif1 (nodes[28], nodes[577],  nodes[639]);
    tranif1 (nodes[364], nodes[738],  nodes[639]);
    tranif1 (nodes[1513], nodes[463],  nodes[639]);
    tranif1 (nodes[558], nodes[1094],  nodes[1630]);
    tranif1 (nodes[1712], nodes[558],  nodes[264]);
    tranif1 (nodes[558], nodes[261],  nodes[461]);
    tranif1 (nodes[558], nodes[726],  nodes[461]);
    tranif1 (nodes[1077], nodes[380],  nodes[879]);
    tranif1 (nodes[558], nodes[238],  nodes[1713]);
    tranif1 (nodes[1354], nodes[623],  nodes[1628]);
    tranif1 (nodes[713], nodes[558],  nodes[907]);
    tranif1 (nodes[1282], nodes[1022],  nodes[414]);
    tranif1 (nodes[1139], nodes[413],  nodes[414]);
    tranif1 (nodes[684], nodes[1359],  nodes[414]);
    tranif1 (nodes[655], nodes[1242],  nodes[414]);
    tranif1 (nodes[1630], nodes[622],  nodes[414]);
    tranif1 (nodes[900], nodes[1437],  nodes[414]);
    tranif1 (nodes[377], nodes[121],  nodes[414]);
    tranif1 (nodes[1185], nodes[558],  nodes[248]);
    tranif1 (nodes[744], nodes[558],  nodes[1108]);
    tranif1 (nodes[558], nodes[140],  nodes[1271]);
    tranif1 (nodes[312], nodes[558],  nodes[159]);
    tranif1 (nodes[1287], nodes[1637],  nodes[129]);
    tranif1 (nodes[1659], nodes[558],  nodes[499]);
    tranif1 (nodes[743], nodes[558],  nodes[499]);
    tranif1 (nodes[558], nodes[252],  nodes[950]);
    tranif1 (nodes[618], nodes[558],  nodes[1029]);
    tranif1 (nodes[695], nodes[1341],  nodes[943]);
    tranif1 (nodes[657], nodes[1237],  nodes[475]);
    tranif1 (nodes[1001], nodes[1435],  nodes[874]);
    tranif1 (nodes[558], nodes[1340],  nodes[642]);
    tranif1 (nodes[558], nodes[1340],  nodes[642]);
    tranif1 (nodes[558], nodes[1340],  nodes[642]);
    tranif1 (nodes[558], nodes[1340],  nodes[642]);
    tranif1 (nodes[558], nodes[152],  nodes[1002]);
    tranif1 (nodes[1407], nodes[558],  nodes[572]);
    tranif1 (nodes[334], nodes[1078],  nodes[943]);
    tranif1 (nodes[657], nodes[451],  nodes[1479]);
    tranif1 (nodes[657], nodes[451],  nodes[1479]);
    tranif1 (nodes[657], nodes[451],  nodes[1479]);
    tranif1 (nodes[451], nodes[657],  nodes[1479]);
    tranif1 (nodes[657], nodes[451],  nodes[1479]);
    tranif1 (nodes[1521], nodes[558],  nodes[1648]);
    tranif1 (nodes[558], nodes[14],  nodes[323]);
    tranif1 (nodes[593], nodes[558],  nodes[355]);
    tranif1 (nodes[1700], nodes[657],  nodes[355]);
    tranif1 (nodes[558], nodes[814],  nodes[392]);
    tranif1 (nodes[558], nodes[557],  nodes[392]);
    tranif1 (nodes[558], nodes[82],  nodes[794]);
    tranif1 (nodes[558], nodes[82],  nodes[794]);
    tranif1 (nodes[82], nodes[558],  nodes[794]);
    tranif1 (nodes[82], nodes[558],  nodes[794]);
    tranif1 (nodes[558], nodes[82],  nodes[794]);
    tranif1 (nodes[558], nodes[82],  nodes[794]);
    tranif1 (nodes[558], nodes[82],  nodes[794]);
    tranif1 (nodes[1436], nodes[1155],  nodes[943]);
    tranif1 (nodes[610], nodes[696],  nodes[943]);
    tranif1 (nodes[558], nodes[811],  nodes[1146]);
    tranif1 (nodes[558], nodes[1440],  nodes[248]);
    tranif1 (nodes[936], nodes[558],  nodes[841]);
    tranif1 (nodes[558], nodes[1501],  nodes[63]);
    tranif1 (nodes[558], nodes[23],  nodes[63]);
    tranif1 (nodes[558], nodes[801],  nodes[1247]);
    tranif1 (nodes[558], nodes[1230],  nodes[43]);
    tranif1 (nodes[558], nodes[570],  nodes[122]);
    tranif1 (nodes[558], nodes[1313],  nodes[649]);
    tranif1 (nodes[558], nodes[640],  nodes[649]);
    tranif1 (nodes[558], nodes[452],  nodes[1332]);
    tranif1 (nodes[558], nodes[1691],  nodes[1332]);
    tranif1 (nodes[558], nodes[1196],  nodes[934]);
    tranif1 (nodes[1585], nodes[558],  nodes[943]);
    tranif1 (nodes[1518], nodes[558],  nodes[1270]);
    tranif1 (nodes[657], nodes[898],  nodes[1270]);
    tranif1 (nodes[558], nodes[432],  nodes[1188]);
    tranif1 (nodes[558], nodes[432],  nodes[1188]);
    tranif1 (nodes[714], nodes[558],  nodes[906]);
    tranif1 (nodes[214], nodes[558],  nodes[906]);
    tranif1 (nodes[578], nodes[558],  nodes[1017]);
    tranif1 (nodes[558], nodes[462],  nodes[1338]);
    tranif1 (nodes[558], nodes[1350],  nodes[1382]);
    tranif1 (nodes[1591], nodes[657],  nodes[7]);
    tranif1 (nodes[1591], nodes[657],  nodes[7]);
    tranif1 (nodes[1591], nodes[657],  nodes[7]);
    tranif1 (nodes[1526], nodes[558],  nodes[680]);
    tranif1 (nodes[760], nodes[629],  nodes[943]);
    tranif1 (nodes[1427], nodes[558],  nodes[967]);
    tranif1 (nodes[558], nodes[852],  nodes[1001]);
    tranif1 (nodes[558], nodes[852],  nodes[1001]);
    tranif1 (nodes[558], nodes[211],  nodes[138]);
    tranif1 (nodes[558], nodes[211],  nodes[138]);
    tranif1 (nodes[558], nodes[211],  nodes[138]);
    tranif1 (nodes[558], nodes[211],  nodes[138]);
    tranif1 (nodes[1027], nodes[1649],  nodes[943]);
    tranif1 (nodes[187], nodes[558],  nodes[926]);
    tranif1 (nodes[604], nodes[1118],  nodes[638]);
    tranif1 (nodes[558], nodes[396],  nodes[1358]);
    tranif1 (nodes[435], nodes[657],  nodes[634]);
    tranif1 (nodes[435], nodes[657],  nodes[634]);
    tranif1 (nodes[435], nodes[657],  nodes[634]);
    tranif1 (nodes[435], nodes[657],  nodes[634]);
    tranif1 (nodes[657], nodes[435],  nodes[634]);
    tranif1 (nodes[1568], nodes[1099],  nodes[1542]);
    tranif1 (nodes[1498], nodes[1184],  nodes[1253]);
    tranif1 (nodes[558], nodes[903],  nodes[1253]);
    tranif1 (nodes[1471], nodes[558],  nodes[827]);
    tranif1 (nodes[558], nodes[392],  nodes[386]);
    tranif1 (nodes[558], nodes[1704],  nodes[386]);
    tranif1 (nodes[1565], nodes[700],  nodes[943]);
    tranif1 (nodes[558], nodes[1166],  nodes[329]);
    tranif1 (nodes[558], nodes[1704],  nodes[329]);
    tranif1 (nodes[558], nodes[1107],  nodes[492]);
    tranif1 (nodes[558], nodes[1005],  nodes[1072]);
    tranif1 (nodes[1005], nodes[558],  nodes[1072]);
    tranif1 (nodes[558], nodes[1005],  nodes[1072]);
    tranif1 (nodes[1005], nodes[558],  nodes[1072]);
    tranif1 (nodes[558], nodes[1005],  nodes[1072]);
    tranif1 (nodes[1005], nodes[558],  nodes[1072]);
    tranif1 (nodes[558], nodes[1005],  nodes[1072]);
    tranif1 (nodes[1005], nodes[558],  nodes[1072]);
    tranif1 (nodes[547], nodes[486],  nodes[1571]);
    tranif1 (nodes[558], nodes[817],  nodes[1571]);
    tranif1 (nodes[657], nodes[230],  nodes[826]);
    tranif1 (nodes[1716], nodes[558],  nodes[218]);
    tranif1 (nodes[688], nodes[1594],  nodes[943]);
    tranif1 (nodes[67], nodes[558],  nodes[1395]);
    tranif1 (nodes[558], nodes[67],  nodes[1395]);
    tranif1 (nodes[1111], nodes[941],  nodes[215]);
    tranif1 (nodes[250], nodes[155],  nodes[59]);
    tranif1 (nodes[669], nodes[558],  nodes[1504]);
    tranif1 (nodes[282], nodes[558],  nodes[6]);
    tranif1 (nodes[657], nodes[874],  nodes[6]);
    tranif1 (nodes[1037], nodes[1280],  nodes[145]);
    tranif1 (nodes[558], nodes[35],  nodes[43]);
    tranif1 (nodes[583], nodes[558],  nodes[991]);
    tranif1 (nodes[558], nodes[730],  nodes[448]);
    tranif1 (nodes[1567], nodes[558],  nodes[678]);
    tranif1 (nodes[1319], nodes[361],  nodes[943]);
    tranif1 (nodes[93], nodes[758],  nodes[943]);
    tranif1 (nodes[558], nodes[1152],  nodes[951]);
    tranif1 (nodes[657], nodes[642],  nodes[951]);
    tranif1 (nodes[657], nodes[1287],  nodes[943]);
    tranif1 (nodes[752], nodes[1190],  nodes[943]);
    tranif1 (nodes[657], nodes[892],  nodes[943]);
    tranif1 (nodes[558], nodes[1130],  nodes[1258]);
    tranif1 (nodes[586], nodes[558],  nodes[1619]);
    tranif1 (nodes[558], nodes[356],  nodes[923]);
    tranif1 (nodes[558], nodes[1334],  nodes[923]);
    tranif1 (nodes[558], nodes[810],  nodes[923]);
    

    supply0 gnd;
    supply1 vcc;
    assign nodes[558] = 1'b0;
    assign nodes[657] = 1'b1;


    assign nodes[159] = reset,
           nodes[89] = ready,
           nodes[1171] = clock0,
           clock1 = nodes[1163],
           clock2 = nodes[421],
           nodes[103] = irq, 
           nodes[1297] = nmi,
           nodes[1672] = so;
     //      sync   =  nodes[];

     assign readNotWrite = nodes[1156] ;
     assign address = {
         nodes[195], 
         nodes[672], 
         nodes[349], 
         nodes[1237], 
         nodes[399], 
         nodes[1443], 
         nodes[148], 
         nodes[230], 
         nodes[1493], 
         nodes[887], 
         nodes[736], 
         nodes[435], 
         nodes[211], 
         nodes[1340], 
         nodes[451], 
         nodes[268]
         
     };

     assign data = {
         nodes[1349], 
         nodes[1591], 
         nodes[175], 
         nodes[1393], 
         nodes[650], 
         nodes[945], 
         nodes[82], 
         nodes[1005]
         
     };

endmodule
