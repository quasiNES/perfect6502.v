module Perfect6502 ( 
    input  reset,
    input  ready,
    input  clock0,
    output clock1,
    output clock2,
    input irq,
    input nmi,
    input so,
    output sync,
    output readNotWrite,
    output [15:0] address,
    inout [7:0] data
);

    wire [3999:0] nodes;

    nmos (nodes[217], nodes[558],  nodes[357]);
    nmos (nodes[349], nodes[657],  nodes[1608]);
    nmos (nodes[1146], nodes[558],  nodes[412]);
    nmos (nodes[943], nodes[558],  nodes[558]);
    nmos (nodes[657], nodes[230],  nodes[826]);
    nmos (nodes[1319], nodes[558],  nodes[82]);
    nmos (nodes[1514], nodes[289],  nodes[821]);
    nmos (nodes[1171], nodes[558],  nodes[558]);
    nmos (nodes[1199], nodes[558],  nodes[945]);
    nmos (nodes[1548], nodes[524],  nodes[710]);
    nmos (nodes[220], nodes[558],  nodes[190]);
    nmos (nodes[657], nodes[1247],  nodes[38]);
    nmos (nodes[558], nodes[189],  nodes[1248]);
    nmos (nodes[155], nodes[558],  nodes[1248]);
    nmos (nodes[346], nodes[558],  nodes[943]);
    nmos (nodes[657], nodes[148],  nodes[1140]);
    nmos (nodes[558], nodes[508],  nodes[1540]);
    nmos (nodes[1082], nodes[32],  nodes[710]);
    nmos (nodes[212], nodes[1451],  nodes[710]);
    nmos (nodes[534], nodes[558],  nodes[1247]);
    nmos (nodes[272], nodes[1162],  nodes[943]);
    nmos (nodes[418], nodes[983],  nodes[943]);
    nmos (nodes[468], nodes[1615],  nodes[248]);
    nmos (nodes[395], nodes[472],  nodes[248]);
    nmos (nodes[348], nodes[1495],  nodes[710]);
    nmos (nodes[558], nodes[1100],  nodes[1096]);
    nmos (nodes[1660], nodes[558],  nodes[1096]);
    nmos (nodes[657], nodes[855],  nodes[1096]);
    nmos (nodes[744], nodes[558],  nodes[1503]);
    nmos (nodes[558], nodes[1616],  nodes[44]);
    nmos (nodes[375], nodes[651],  nodes[78]);
    nmos (nodes[65], nodes[558],  nodes[78]);
    nmos (nodes[1378], nodes[928],  nodes[710]);
    nmos (nodes[74], nodes[1309],  nodes[710]);
    nmos (nodes[115], nodes[518],  nodes[943]);
    nmos (nodes[31], nodes[558],  nodes[32]);
    nmos (nodes[657], nodes[1405],  nodes[943]);
    nmos (nodes[1603], nodes[973],  nodes[943]);
    nmos (nodes[558], nodes[510],  nodes[347]);
    nmos (nodes[883], nodes[1667],  nodes[710]);
    nmos (nodes[558], nodes[1456],  nodes[706]);
    nmos (nodes[558], nodes[307],  nodes[1174]);
    nmos (nodes[409], nodes[558],  nodes[1622]);
    nmos (nodes[558], nodes[25],  nodes[192]);
    nmos (nodes[606], nodes[558],  nodes[1490]);
    nmos (nodes[767], nodes[1148],  nodes[943]);
    nmos (nodes[1248], nodes[1150],  nodes[549]);
    nmos (nodes[1332], nodes[1287],  nodes[549]);
    nmos (nodes[1188], nodes[1680],  nodes[549]);
    nmos (nodes[1405], nodes[1142],  nodes[549]);
    nmos (nodes[558], nodes[794],  nodes[353]);
    nmos (nodes[558], nodes[794],  nodes[353]);
    nmos (nodes[1700], nodes[558],  nodes[593]);
    nmos (nodes[54], nodes[1167],  nodes[549]);
    nmos (nodes[1362], nodes[613],  nodes[600]);
    nmos (nodes[166], nodes[530],  nodes[549]);
    nmos (nodes[1336], nodes[1627],  nodes[549]);
    nmos (nodes[1400], nodes[558],  nodes[948]);
    nmos (nodes[480], nodes[1092],  nodes[264]);
    nmos (nodes[558], nodes[632],  nodes[1582]);
    nmos (nodes[923], nodes[558],  nodes[584]);
    nmos (nodes[136], nodes[274],  nodes[1003]);
    nmos (nodes[558], nodes[860],  nodes[1003]);
    nmos (nodes[1527], nodes[1347],  nodes[943]);
    nmos (nodes[331], nodes[558],  nodes[68]);
    nmos (nodes[558], nodes[945],  nodes[558]);
    nmos (nodes[1495], nodes[1644],  nodes[1457]);
    nmos (nodes[558], nodes[1066],  nodes[1485]);
    nmos (nodes[1066], nodes[558],  nodes[1485]);
    nmos (nodes[558], nodes[1066],  nodes[1485]);
    nmos (nodes[1622], nodes[558],  nodes[1077]);
    nmos (nodes[558], nodes[667],  nodes[1077]);
    nmos (nodes[1336], nodes[115],  nodes[325]);
    nmos (nodes[785], nodes[920],  nodes[710]);
    nmos (nodes[558], nodes[748],  nodes[1318]);
    nmos (nodes[657], nodes[304],  nodes[362]);
    nmos (nodes[657], nodes[421],  nodes[127]);
    nmos (nodes[1405], nodes[989],  nodes[325]);
    nmos (nodes[790], nodes[558],  nodes[53]);
    nmos (nodes[1068], nodes[558],  nodes[763]);
    nmos (nodes[147], nodes[558],  nodes[1088]);
    nmos (nodes[1463], nodes[558],  nodes[1088]);
    nmos (nodes[493], nodes[1370],  nodes[1042]);
    nmos (nodes[1421], nodes[1473],  nodes[1042]);
    nmos (nodes[443], nodes[513],  nodes[943]);
    nmos (nodes[1646], nodes[1673],  nodes[943]);
    nmos (nodes[1516], nodes[490],  nodes[943]);
    nmos (nodes[558], nodes[856],  nodes[311]);
    nmos (nodes[558], nodes[835],  nodes[311]);
    nmos (nodes[1158], nodes[558],  nodes[783]);
    nmos (nodes[1704], nodes[558],  nodes[783]);
    nmos (nodes[1253], nodes[558],  nodes[783]);
    nmos (nodes[558], nodes[230],  nodes[381]);
    nmos (nodes[558], nodes[230],  nodes[381]);
    nmos (nodes[558], nodes[230],  nodes[381]);
    nmos (nodes[230], nodes[558],  nodes[381]);
    nmos (nodes[558], nodes[230],  nodes[381]);
    nmos (nodes[230], nodes[558],  nodes[381]);
    nmos (nodes[558], nodes[230],  nodes[381]);
    nmos (nodes[1343], nodes[558],  nodes[152]);
    nmos (nodes[558], nodes[371],  nodes[555]);
    nmos (nodes[207], nodes[558],  nodes[810]);
    nmos (nodes[558], nodes[501],  nodes[819]);
    nmos (nodes[558], nodes[1138],  nodes[1148]);
    nmos (nodes[672], nodes[657],  nodes[963]);
    nmos (nodes[558], nodes[202],  nodes[967]);
    nmos (nodes[558], nodes[972],  nodes[1691]);
    nmos (nodes[558], nodes[1563],  nodes[1342]);
    nmos (nodes[558], nodes[844],  nodes[786]);
    nmos (nodes[1296], nodes[657],  nodes[422]);
    nmos (nodes[558], nodes[1346],  nodes[422]);
    nmos (nodes[558], nodes[359],  nodes[422]);
    nmos (nodes[558], nodes[1680],  nodes[984]);
    nmos (nodes[365], nodes[558],  nodes[1410]);
    nmos (nodes[1145], nodes[558],  nodes[403]);
    nmos (nodes[558], nodes[746],  nodes[527]);
    nmos (nodes[1372], nodes[972],  nodes[1610]);
    nmos (nodes[1497], nodes[653],  nodes[710]);
    nmos (nodes[558], nodes[489],  nodes[429]);
    nmos (nodes[10], nodes[558],  nodes[467]);
    nmos (nodes[558], nodes[692],  nodes[460]);
    nmos (nodes[1647], nodes[558],  nodes[536]);
    nmos (nodes[558], nodes[1358],  nodes[917]);
    nmos (nodes[514], nodes[429],  nodes[821]);
    nmos (nodes[1268], nodes[558],  nodes[744]);
    nmos (nodes[1570], nodes[430],  nodes[710]);
    nmos (nodes[393], nodes[1179],  nodes[943]);
    nmos (nodes[1188], nodes[998],  nodes[1700]);
    nmos (nodes[1287], nodes[1389],  nodes[1700]);
    nmos (nodes[1462], nodes[558],  nodes[1369]);
    nmos (nodes[438], nodes[657],  nodes[1369]);
    nmos (nodes[816], nodes[558],  nodes[925]);
    nmos (nodes[1001], nodes[721],  nodes[1700]);
    nmos (nodes[1336], nodes[618],  nodes[1700]);
    nmos (nodes[558], nodes[1043],  nodes[818]);
    nmos (nodes[414], nodes[657],  nodes[818]);
    nmos (nodes[1405], nodes[3],  nodes[1700]);
    nmos (nodes[558], nodes[1426],  nodes[270]);
    nmos (nodes[1559], nodes[477],  nodes[1678]);
    nmos (nodes[1632], nodes[558],  nodes[1678]);
    nmos (nodes[1083], nodes[1590],  nodes[710]);
    nmos (nodes[1017], nodes[558],  nodes[589]);
    nmos (nodes[1066], nodes[1424],  nodes[710]);
    nmos (nodes[558], nodes[1455],  nodes[1420]);
    nmos (nodes[558], nodes[397],  nodes[1420]);
    nmos (nodes[558], nodes[789],  nodes[493]);
    nmos (nodes[558], nodes[884],  nodes[640]);
    nmos (nodes[624], nodes[558],  nodes[1108]);
    nmos (nodes[75], nodes[558],  nodes[154]);
    nmos (nodes[129], nodes[657],  nodes[154]);
    nmos (nodes[605], nodes[558],  nodes[787]);
    nmos (nodes[325], nodes[558],  nodes[1247]);
    nmos (nodes[558], nodes[604],  nodes[1582]);
    nmos (nodes[558], nodes[1010],  nodes[1670]);
    nmos (nodes[657], nodes[82],  nodes[798]);
    nmos (nodes[657], nodes[82],  nodes[798]);
    nmos (nodes[558], nodes[1264],  nodes[453]);
    nmos (nodes[558], nodes[567],  nodes[28]);
    nmos (nodes[1548], nodes[558],  nodes[121]);
    nmos (nodes[558], nodes[1225],  nodes[285]);
    nmos (nodes[70], nodes[558],  nodes[1134]);
    nmos (nodes[558], nodes[1366],  nodes[706]);
    nmos (nodes[558], nodes[952],  nodes[272]);
    nmos (nodes[558], nodes[426],  nodes[715]);
    nmos (nodes[558], nodes[914],  nodes[715]);
    nmos (nodes[739], nodes[711],  nodes[761]);
    nmos (nodes[399], nodes[657],  nodes[1296]);
    nmos (nodes[373], nodes[657],  nodes[1453]);
    nmos (nodes[264], nodes[558],  nodes[1312]);
    nmos (nodes[812], nodes[558],  nodes[646]);
    nmos (nodes[210], nodes[1513],  nodes[943]);
    nmos (nodes[1706], nodes[1500],  nodes[379]);
    nmos (nodes[1345], nodes[558],  nodes[379]);
    nmos (nodes[1508], nodes[1101],  nodes[813]);
    nmos (nodes[11], nodes[558],  nodes[4]);
    nmos (nodes[558], nodes[1380],  nodes[819]);
    nmos (nodes[657], nodes[214],  nodes[714]);
    nmos (nodes[558], nodes[818],  nodes[43]);
    nmos (nodes[1107], nodes[558],  nodes[1520]);
    nmos (nodes[1130], nodes[558],  nodes[1002]);
    nmos (nodes[805], nodes[779],  nodes[943]);
    nmos (nodes[101], nodes[1141],  nodes[710]);
    nmos (nodes[1308], nodes[408],  nodes[943]);
    nmos (nodes[379], nodes[1480],  nodes[1581]);
    nmos (nodes[191], nodes[558],  nodes[347]);
    nmos (nodes[558], nodes[1116],  nodes[1537]);
    nmos (nodes[1116], nodes[558],  nodes[1537]);
    nmos (nodes[558], nodes[1116],  nodes[1537]);
    nmos (nodes[558], nodes[169],  nodes[1624]);
    nmos (nodes[558], nodes[938],  nodes[408]);
    nmos (nodes[558], nodes[1125],  nodes[1576]);
    nmos (nodes[1394], nodes[1609],  nodes[943]);
    nmos (nodes[558], nodes[453],  nodes[205]);
    nmos (nodes[368], nodes[558],  nodes[309]);
    nmos (nodes[1172], nodes[405],  nodes[1544]);
    nmos (nodes[373], nodes[558],  nodes[1720]);
    nmos (nodes[612], nodes[657],  nodes[1720]);
    nmos (nodes[657], nodes[1076],  nodes[1088]);
    nmos (nodes[773], nodes[558],  nodes[646]);
    nmos (nodes[1141], nodes[558],  nodes[982]);
    nmos (nodes[1203], nodes[558],  nodes[1135]);
    nmos (nodes[1629], nodes[558],  nodes[1135]);
    nmos (nodes[813], nodes[558],  nodes[1258]);
    nmos (nodes[720], nodes[558],  nodes[248]);
    nmos (nodes[1371], nodes[558],  nodes[1045]);
    nmos (nodes[1237], nodes[558],  nodes[999]);
    nmos (nodes[558], nodes[1237],  nodes[999]);
    nmos (nodes[1237], nodes[558],  nodes[999]);
    nmos (nodes[1237], nodes[558],  nodes[999]);
    nmos (nodes[558], nodes[1237],  nodes[999]);
    nmos (nodes[1237], nodes[558],  nodes[999]);
    nmos (nodes[558], nodes[1237],  nodes[999]);
    nmos (nodes[29], nodes[561],  nodes[943]);
    nmos (nodes[876], nodes[558],  nodes[867]);
    nmos (nodes[1717], nodes[558],  nodes[1173]);
    nmos (nodes[558], nodes[206],  nodes[1146]);
    nmos (nodes[1106], nodes[558],  nodes[76]);
    nmos (nodes[1033], nodes[558],  nodes[241]);
    nmos (nodes[1015], nodes[657],  nodes[241]);
    nmos (nodes[886], nodes[975],  nodes[995]);
    nmos (nodes[1371], nodes[558],  nodes[201]);
    nmos (nodes[272], nodes[558],  nodes[273]);
    nmos (nodes[558], nodes[307],  nodes[846]);
    nmos (nodes[541], nodes[1183],  nodes[879]);
    nmos (nodes[380], nodes[558],  nodes[827]);
    nmos (nodes[124], nodes[558],  nodes[1061]);
    nmos (nodes[1403], nodes[332],  nodes[654]);
    nmos (nodes[657], nodes[1108],  nodes[943]);
    nmos (nodes[355], nodes[558],  nodes[621]);
    nmos (nodes[251], nodes[558],  nodes[1035]);
    nmos (nodes[558], nodes[188],  nodes[1606]);
    nmos (nodes[719], nodes[407],  nodes[41]);
    nmos (nodes[87], nodes[52],  nodes[41]);
    nmos (nodes[1424], nodes[1651],  nodes[41]);
    nmos (nodes[1661], nodes[315],  nodes[41]);
    nmos (nodes[1095], nodes[1160],  nodes[41]);
    nmos (nodes[1387], nodes[483],  nodes[41]);
    nmos (nodes[1014], nodes[13],  nodes[41]);
    nmos (nodes[1147], nodes[1539],  nodes[41]);
    nmos (nodes[689], nodes[558],  nodes[370]);
    nmos (nodes[1534], nodes[558],  nodes[805]);
    nmos (nodes[1136], nodes[326],  nodes[943]);
    nmos (nodes[170], nodes[1117],  nodes[943]);
    nmos (nodes[873], nodes[797],  nodes[710]);
    nmos (nodes[1087], nodes[558],  nodes[1382]);
    nmos (nodes[558], nodes[1178],  nodes[960]);
    nmos (nodes[316], nodes[1628],  nodes[977]);
    nmos (nodes[143], nodes[558],  nodes[977]);
    nmos (nodes[166], nodes[1098],  nodes[874]);
    nmos (nodes[1336], nodes[1212],  nodes[874]);
    nmos (nodes[1188], nodes[1532],  nodes[874]);
    nmos (nodes[1702], nodes[1405],  nodes[874]);
    nmos (nodes[1150], nodes[183],  nodes[874]);
    nmos (nodes[1287], nodes[81],  nodes[874]);
    nmos (nodes[558], nodes[802],  nodes[781]);
    nmos (nodes[406], nodes[558],  nodes[1525]);
    nmos (nodes[555], nodes[558],  nodes[1525]);
    nmos (nodes[558], nodes[427],  nodes[647]);
    nmos (nodes[558], nodes[1425],  nodes[1372]);
    nmos (nodes[1648], nodes[242],  nodes[943]);
    nmos (nodes[1674], nodes[931],  nodes[710]);
    nmos (nodes[1450], nodes[1526],  nodes[710]);
    nmos (nodes[558], nodes[638],  nodes[1273]);
    nmos (nodes[154], nodes[558],  nodes[512]);
    nmos (nodes[558], nodes[874],  nodes[1247]);
    nmos (nodes[1448], nodes[558],  nodes[1427]);
    nmos (nodes[1357], nodes[558],  nodes[223]);
    nmos (nodes[1002], nodes[558],  nodes[1219]);
    nmos (nodes[687], nodes[1108],  nodes[1042]);
    nmos (nodes[1477], nodes[604],  nodes[943]);
    nmos (nodes[1082], nodes[367],  nodes[206]);
    nmos (nodes[558], nodes[818],  nodes[265]);
    nmos (nodes[971], nodes[558],  nodes[1575]);
    nmos (nodes[406], nodes[371],  nodes[105]);
    nmos (nodes[555], nodes[558],  nodes[105]);
    nmos (nodes[1323], nodes[558],  nodes[631]);
    nmos (nodes[283], nodes[657],  nodes[631]);
    nmos (nodes[558], nodes[267],  nodes[544]);
    nmos (nodes[558], nodes[616],  nodes[1482]);
    nmos (nodes[1437], nodes[657],  nodes[943]);
    nmos (nodes[1364], nodes[558],  nodes[101]);
    nmos (nodes[844], nodes[558],  nodes[985]);
    nmos (nodes[1151], nodes[558],  nodes[1262]);
    nmos (nodes[1212], nodes[618],  nodes[654]);
    nmos (nodes[1098], nodes[280],  nodes[654]);
    nmos (nodes[1702], nodes[3],  nodes[654]);
    nmos (nodes[1532], nodes[998],  nodes[654]);
    nmos (nodes[81], nodes[1389],  nodes[654]);
    nmos (nodes[183], nodes[694],  nodes[654]);
    nmos (nodes[883], nodes[558],  nodes[315]);
    nmos (nodes[178], nodes[558],  nodes[1307]);
    nmos (nodes[347], nodes[558],  nodes[281]);
    nmos (nodes[558], nodes[553],  nodes[781]);
    nmos (nodes[1235], nodes[558],  nodes[1413]);
    nmos (nodes[1649], nodes[558],  nodes[764]);
    nmos (nodes[1187], nodes[558],  nodes[1212]);
    nmos (nodes[1597], nodes[719],  nodes[710]);
    nmos (nodes[1605], nodes[558],  nodes[1410]);
    nmos (nodes[558], nodes[455],  nodes[279]);
    nmos (nodes[657], nodes[407],  nodes[943]);
    nmos (nodes[558], nodes[1724],  nodes[730]);
    nmos (nodes[175], nodes[558],  nodes[612]);
    nmos (nodes[175], nodes[558],  nodes[612]);
    nmos (nodes[175], nodes[558],  nodes[612]);
    nmos (nodes[175], nodes[558],  nodes[612]);
    nmos (nodes[558], nodes[175],  nodes[612]);
    nmos (nodes[558], nodes[175],  nodes[612]);
    nmos (nodes[175], nodes[558],  nodes[612]);
    nmos (nodes[317], nodes[558],  nodes[445]);
    nmos (nodes[417], nodes[558],  nodes[445]);
    nmos (nodes[417], nodes[558],  nodes[445]);
    nmos (nodes[558], nodes[127],  nodes[710]);
    nmos (nodes[558], nodes[539],  nodes[445]);
    nmos (nodes[539], nodes[558],  nodes[445]);
    nmos (nodes[558], nodes[539],  nodes[445]);
    nmos (nodes[539], nodes[558],  nodes[445]);
    nmos (nodes[539], nodes[558],  nodes[445]);
    nmos (nodes[558], nodes[287],  nodes[768]);
    nmos (nodes[558], nodes[1215],  nodes[1382]);
    nmos (nodes[547], nodes[558],  nodes[1220]);
    nmos (nodes[558], nodes[817],  nodes[1220]);
    nmos (nodes[1242], nodes[1637],  nodes[1015]);
    nmos (nodes[872], nodes[1282],  nodes[1015]);
    nmos (nodes[401], nodes[413],  nodes[1015]);
    nmos (nodes[1464], nodes[558],  nodes[784]);
    nmos (nodes[501], nodes[558],  nodes[67]);
    nmos (nodes[913], nodes[558],  nodes[1699]);
    nmos (nodes[558], nodes[261],  nodes[447]);
    nmos (nodes[558], nodes[388],  nodes[425]);
    nmos (nodes[54], nodes[564],  nodes[801]);
    nmos (nodes[558], nodes[335],  nodes[347]);
    nmos (nodes[1596], nodes[558],  nodes[1602]);
    nmos (nodes[558], nodes[442],  nodes[182]);
    nmos (nodes[798], nodes[657],  nodes[746]);
    nmos (nodes[729], nodes[261],  nodes[943]);
    nmos (nodes[323], nodes[959],  nodes[710]);
    nmos (nodes[1605], nodes[1183],  nodes[710]);
    nmos (nodes[793], nodes[1181],  nodes[1595]);
    nmos (nodes[558], nodes[488],  nodes[1227]);
    nmos (nodes[558], nodes[182],  nodes[0]);
    nmos (nodes[558], nodes[861],  nodes[1452]);
    nmos (nodes[1000], nodes[558],  nodes[575]);
    nmos (nodes[1055], nodes[558],  nodes[1708]);
    nmos (nodes[921], nodes[558],  nodes[1305]);
    nmos (nodes[558], nodes[800],  nodes[525]);
    nmos (nodes[657], nodes[1331],  nodes[525]);
    nmos (nodes[558], nodes[80],  nodes[1130]);
    nmos (nodes[980], nodes[558],  nodes[1381]);
    nmos (nodes[558], nodes[1133],  nodes[328]);
    nmos (nodes[194], nodes[558],  nodes[328]);
    nmos (nodes[558], nodes[451],  nodes[66]);
    nmos (nodes[558], nodes[451],  nodes[66]);
    nmos (nodes[558], nodes[451],  nodes[66]);
    nmos (nodes[558], nodes[451],  nodes[66]);
    nmos (nodes[48], nodes[558],  nodes[943]);
    nmos (nodes[741], nodes[558],  nodes[943]);
    nmos (nodes[558], nodes[600],  nodes[1341]);
    nmos (nodes[300], nodes[558],  nodes[712]);
    nmos (nodes[1224], nodes[558],  nodes[1108]);
    nmos (nodes[1397], nodes[1303],  nodes[335]);
    nmos (nodes[558], nodes[279],  nodes[253]);
    nmos (nodes[558], nodes[1692],  nodes[253]);
    nmos (nodes[943], nodes[657],  nodes[1129]);
    nmos (nodes[558], nodes[906],  nodes[1333]);
    nmos (nodes[558], nodes[82],  nodes[558]);
    nmos (nodes[605], nodes[558],  nodes[1081]);
    nmos (nodes[1198], nodes[558],  nodes[1530]);
    nmos (nodes[248], nodes[657],  nodes[424]);
    nmos (nodes[1178], nodes[558],  nodes[614]);
    nmos (nodes[558], nodes[248],  nodes[198]);
    nmos (nodes[558], nodes[424],  nodes[198]);
    nmos (nodes[1604], nodes[1717],  nodes[335]);
    nmos (nodes[977], nodes[413],  nodes[437]);
    nmos (nodes[1054], nodes[558],  nodes[926]);
    nmos (nodes[1150], nodes[694],  nodes[1700]);
    nmos (nodes[349], nodes[558],  nodes[869]);
    nmos (nodes[349], nodes[558],  nodes[869]);
    nmos (nodes[558], nodes[349],  nodes[869]);
    nmos (nodes[349], nodes[558],  nodes[869]);
    nmos (nodes[558], nodes[349],  nodes[869]);
    nmos (nodes[558], nodes[349],  nodes[869]);
    nmos (nodes[558], nodes[349],  nodes[869]);
    nmos (nodes[1393], nodes[657],  nodes[1076]);
    nmos (nodes[1393], nodes[657],  nodes[1076]);
    nmos (nodes[641], nodes[558],  nodes[1611]);
    nmos (nodes[166], nodes[280],  nodes[1700]);
    nmos (nodes[544], nodes[558],  nodes[244]);
    nmos (nodes[939], nodes[757],  nodes[1144]);
    nmos (nodes[428], nodes[1456],  nodes[248]);
    nmos (nodes[1091], nodes[12],  nodes[248]);
    nmos (nodes[16], nodes[558],  nodes[248]);
    nmos (nodes[558], nodes[213],  nodes[82]);
    nmos (nodes[686], nodes[558],  nodes[170]);
    nmos (nodes[280], nodes[558],  nodes[601]);
    nmos (nodes[162], nodes[1654],  nodes[943]);
    nmos (nodes[1062], nodes[705],  nodes[821]);
    nmos (nodes[558], nodes[6],  nodes[521]);
    nmos (nodes[417], nodes[657],  nodes[317]);
    nmos (nodes[52], nodes[558],  nodes[203]);
    nmos (nodes[1076], nodes[558],  nodes[353]);
    nmos (nodes[1076], nodes[558],  nodes[353]);
    nmos (nodes[1463], nodes[558],  nodes[353]);
    nmos (nodes[845], nodes[1553],  nodes[710]);
    nmos (nodes[558], nodes[1358],  nodes[1109]);
    nmos (nodes[1281], nodes[558],  nodes[650]);
    nmos (nodes[500], nodes[558],  nodes[427]);
    nmos (nodes[1314], nodes[112],  nodes[427]);
    nmos (nodes[462], nodes[878],  nodes[943]);
    nmos (nodes[558], nodes[807],  nodes[330]);
    nmos (nodes[1716], nodes[558],  nodes[1258]);
    nmos (nodes[315], nodes[584],  nodes[48]);
    nmos (nodes[1651], nodes[502],  nodes[48]);
    nmos (nodes[483], nodes[49],  nodes[48]);
    nmos (nodes[1160], nodes[948],  nodes[48]);
    nmos (nodes[1539], nodes[205],  nodes[48]);
    nmos (nodes[13], nodes[1551],  nodes[48]);
    nmos (nodes[657], nodes[1336],  nodes[943]);
    nmos (nodes[1029], nodes[1187],  nodes[943]);
    nmos (nodes[1383], nodes[558],  nodes[1503]);
    nmos (nodes[92], nodes[1667],  nodes[821]);
    nmos (nodes[1683], nodes[1090],  nodes[943]);
    nmos (nodes[1018], nodes[558],  nodes[762]);
    nmos (nodes[558], nodes[421],  nodes[135]);
    nmos (nodes[558], nodes[421],  nodes[135]);
    nmos (nodes[421], nodes[558],  nodes[135]);
    nmos (nodes[558], nodes[421],  nodes[135]);
    nmos (nodes[657], nodes[1160],  nodes[943]);
    nmos (nodes[657], nodes[1630],  nodes[943]);
    nmos (nodes[1012], nodes[366],  nodes[440]);
    nmos (nodes[558], nodes[1143],  nodes[668]);
    nmos (nodes[558], nodes[21],  nodes[1162]);
    nmos (nodes[15], nodes[474],  nodes[943]);
    nmos (nodes[54], nodes[1169],  nodes[1263]);
    nmos (nodes[1035], nodes[558],  nodes[962]);
    nmos (nodes[558], nodes[963],  nodes[1523]);
    nmos (nodes[657], nodes[635],  nodes[1523]);
    nmos (nodes[558], nodes[1413],  nodes[1260]);
    nmos (nodes[1235], nodes[657],  nodes[1260]);
    nmos (nodes[130], nodes[558],  nodes[220]);
    nmos (nodes[657], nodes[639],  nodes[220]);
    nmos (nodes[102], nodes[558],  nodes[400]);
    nmos (nodes[1696], nodes[657],  nodes[400]);
    nmos (nodes[1696], nodes[558],  nodes[834]);
    nmos (nodes[400], nodes[558],  nodes[834]);
    nmos (nodes[558], nodes[1561],  nodes[777]);
    nmos (nodes[558], nodes[656],  nodes[604]);
    nmos (nodes[657], nodes[1443],  nodes[1545]);
    nmos (nodes[1012], nodes[558],  nodes[1246]);
    nmos (nodes[949], nodes[558],  nodes[1334]);
    nmos (nodes[1406], nodes[558],  nodes[1334]);
    nmos (nodes[1108], nodes[977],  nodes[859]);
    nmos (nodes[187], nodes[402],  nodes[710]);
    nmos (nodes[1129], nodes[558],  nodes[358]);
    nmos (nodes[1129], nodes[558],  nodes[358]);
    nmos (nodes[1113], nodes[1717],  nodes[943]);
    nmos (nodes[1001], nodes[871],  nodes[1263]);
    nmos (nodes[52], nodes[657],  nodes[943]);
    nmos (nodes[498], nodes[568],  nodes[943]);
    nmos (nodes[558], nodes[138],  nodes[1250]);
    nmos (nodes[558], nodes[990],  nodes[1250]);
    nmos (nodes[657], nodes[1041],  nodes[1250]);
    nmos (nodes[1214], nodes[558],  nodes[1011]);
    nmos (nodes[182], nodes[558],  nodes[1655]);
    nmos (nodes[558], nodes[1356],  nodes[1136]);
    nmos (nodes[558], nodes[909],  nodes[378]);
    nmos (nodes[558], nodes[71],  nodes[35]);
    nmos (nodes[657], nodes[654],  nodes[35]);
    nmos (nodes[558], nodes[1180],  nodes[554]);
    nmos (nodes[964], nodes[558],  nodes[554]);
    nmos (nodes[558], nodes[1304],  nodes[787]);
    nmos (nodes[558], nodes[1347],  nodes[967]);
    nmos (nodes[104], nodes[558],  nodes[967]);
    nmos (nodes[343], nodes[571],  nodes[710]);
    nmos (nodes[1061], nodes[207],  nodes[943]);
    nmos (nodes[1004], nodes[473],  nodes[980]);
    nmos (nodes[958], nodes[558],  nodes[89]);
    nmos (nodes[672], nodes[657],  nodes[963]);
    nmos (nodes[558], nodes[863],  nodes[1240]);
    nmos (nodes[333], nodes[164],  nodes[943]);
    nmos (nodes[1197], nodes[558],  nodes[174]);
    nmos (nodes[1170], nodes[558],  nodes[781]);
    nmos (nodes[657], nodes[1417],  nodes[670]);
    nmos (nodes[1443], nodes[558],  nodes[994]);
    nmos (nodes[558], nodes[1443],  nodes[994]);
    nmos (nodes[1443], nodes[558],  nodes[994]);
    nmos (nodes[1443], nodes[558],  nodes[994]);
    nmos (nodes[558], nodes[1443],  nodes[994]);
    nmos (nodes[1443], nodes[558],  nodes[994]);
    nmos (nodes[558], nodes[1443],  nodes[994]);
    nmos (nodes[518], nodes[558],  nodes[1439]);
    nmos (nodes[721], nodes[1435],  nodes[654]);
    nmos (nodes[880], nodes[558],  nodes[13]);
    nmos (nodes[558], nodes[747],  nodes[670]);
    nmos (nodes[558], nodes[1480],  nodes[1472]);
    nmos (nodes[558], nodes[1294],  nodes[1587]);
    nmos (nodes[1083], nodes[558],  nodes[1587]);
    nmos (nodes[942], nodes[1285],  nodes[1628]);
    nmos (nodes[877], nodes[558],  nodes[506]);
    nmos (nodes[1642], nodes[1278],  nodes[824]);
    nmos (nodes[1084], nodes[722],  nodes[59]);
    nmos (nodes[558], nodes[1347],  nodes[1396]);
    nmos (nodes[634], nodes[558],  nodes[1676]);
    nmos (nodes[657], nodes[86],  nodes[1676]);
    nmos (nodes[310], nodes[194],  nodes[943]);
    nmos (nodes[558], nodes[1092],  nodes[118]);
    nmos (nodes[572], nodes[558],  nodes[1176]);
    nmos (nodes[558], nodes[61],  nodes[1336]);
    nmos (nodes[558], nodes[268],  nodes[1100]);
    nmos (nodes[558], nodes[268],  nodes[1100]);
    nmos (nodes[558], nodes[268],  nodes[1100]);
    nmos (nodes[383], nodes[558],  nodes[712]);
    nmos (nodes[558], nodes[1560],  nodes[1337]);
    nmos (nodes[3], nodes[558],  nodes[1603]);
    nmos (nodes[754], nodes[1422],  nodes[443]);
    nmos (nodes[755], nodes[558],  nodes[443]);
    nmos (nodes[601], nodes[496],  nodes[943]);
    nmos (nodes[558], nodes[225],  nodes[1223]);
    nmos (nodes[859], nodes[657],  nodes[1223]);
    nmos (nodes[558], nodes[895],  nodes[337]);
    nmos (nodes[1222], nodes[558],  nodes[1225]);
    nmos (nodes[870], nodes[87],  nodes[710]);
    nmos (nodes[1414], nodes[684],  nodes[1015]);
    nmos (nodes[606], nodes[1437],  nodes[1015]);
    nmos (nodes[459], nodes[844],  nodes[943]);
    nmos (nodes[558], nodes[568],  nodes[175]);
    nmos (nodes[558], nodes[916],  nodes[1517]);
    nmos (nodes[1299], nodes[765],  nodes[1015]);
    nmos (nodes[314], nodes[1630],  nodes[1015]);
    nmos (nodes[331], nodes[121],  nodes[1015]);
    nmos (nodes[57], nodes[1402],  nodes[293]);
    nmos (nodes[356], nodes[207],  nodes[293]);
    nmos (nodes[558], nodes[810],  nodes[293]);
    nmos (nodes[1106], nodes[734],  nodes[335]);
    nmos (nodes[558], nodes[330],  nodes[807]);
    nmos (nodes[558], nodes[1041],  nodes[990]);
    nmos (nodes[657], nodes[138],  nodes[990]);
    nmos (nodes[1575], nodes[558],  nodes[1357]);
    nmos (nodes[1475], nodes[558],  nodes[1097]);
    nmos (nodes[1691], nodes[740],  nodes[59]);
    nmos (nodes[29], nodes[51],  nodes[787]);
    nmos (nodes[203], nodes[558],  nodes[1635]);
    nmos (nodes[237], nodes[1641],  nodes[710]);
    nmos (nodes[409], nodes[724],  nodes[710]);
    nmos (nodes[845], nodes[1426],  nodes[1662]);
    nmos (nodes[80], nodes[558],  nodes[267]);
    nmos (nodes[916], nodes[387],  nodes[206]);
    nmos (nodes[1071], nodes[649],  nodes[59]);
    nmos (nodes[1572], nodes[22],  nodes[505]);
    nmos (nodes[193], nodes[558],  nodes[505]);
    nmos (nodes[495], nodes[1071],  nodes[943]);
    nmos (nodes[558], nodes[1130],  nodes[1109]);
    nmos (nodes[558], nodes[1163],  nodes[1417]);
    nmos (nodes[1163], nodes[558],  nodes[1417]);
    nmos (nodes[558], nodes[1163],  nodes[1417]);
    nmos (nodes[1163], nodes[558],  nodes[1417]);
    nmos (nodes[558], nodes[1163],  nodes[1417]);
    nmos (nodes[116], nodes[718],  nodes[943]);
    nmos (nodes[558], nodes[165],  nodes[1236]);
    nmos (nodes[345], nodes[1584],  nodes[8]);
    nmos (nodes[37], nodes[558],  nodes[1634]);
    nmos (nodes[224], nodes[558],  nodes[1634]);
    nmos (nodes[558], nodes[176],  nodes[10]);
    nmos (nodes[558], nodes[628],  nodes[55]);
    nmos (nodes[1616], nodes[299],  nodes[1614]);
    nmos (nodes[335], nodes[558],  nodes[925]);
    nmos (nodes[1697], nodes[558],  nodes[664]);
    nmos (nodes[1134], nodes[558],  nodes[1465]);
    nmos (nodes[558], nodes[122],  nodes[1459]);
    nmos (nodes[558], nodes[1030],  nodes[1459]);
    nmos (nodes[1305], nodes[558],  nodes[772]);
    nmos (nodes[921], nodes[657],  nodes[772]);
    nmos (nodes[496], nodes[558],  nodes[1098]);
    nmos (nodes[558], nodes[481],  nodes[1079]);
    nmos (nodes[558], nodes[534],  nodes[943]);
    nmos (nodes[558], nodes[625],  nodes[459]);
    nmos (nodes[558], nodes[830],  nodes[43]);
    nmos (nodes[558], nodes[103],  nodes[558]);
    nmos (nodes[580], nodes[566],  nodes[755]);
    nmos (nodes[657], nodes[520],  nodes[1634]);
    nmos (nodes[17], nodes[558],  nodes[732]);
    nmos (nodes[1536], nodes[558],  nodes[732]);
    nmos (nodes[1679], nodes[248],  nodes[710]);
    nmos (nodes[1215], nodes[223],  nodes[710]);
    nmos (nodes[558], nodes[1327],  nodes[748]);
    nmos (nodes[511], nodes[558],  nodes[1078]);
    nmos (nodes[719], nodes[1108],  nodes[863]);
    nmos (nodes[87], nodes[991],  nodes[863]);
    nmos (nodes[1424], nodes[1473],  nodes[863]);
    nmos (nodes[1661], nodes[1302],  nodes[863]);
    nmos (nodes[1095], nodes[892],  nodes[863]);
    nmos (nodes[1387], nodes[1503],  nodes[863]);
    nmos (nodes[1014], nodes[833],  nodes[863]);
    nmos (nodes[1147], nodes[493],  nodes[863]);
    nmos (nodes[558], nodes[1368],  nodes[1374]);
    nmos (nodes[1493], nodes[657],  nodes[322]);
    nmos (nodes[657], nodes[1493],  nodes[322]);
    nmos (nodes[657], nodes[1493],  nodes[322]);
    nmos (nodes[657], nodes[1493],  nodes[322]);
    nmos (nodes[1233], nodes[558],  nodes[1536]);
    nmos (nodes[286], nodes[558],  nodes[1536]);
    nmos (nodes[382], nodes[558],  nodes[1536]);
    nmos (nodes[1173], nodes[558],  nodes[1536]);
    nmos (nodes[1543], nodes[558],  nodes[1536]);
    nmos (nodes[76], nodes[558],  nodes[1536]);
    nmos (nodes[558], nodes[1658],  nodes[1536]);
    nmos (nodes[558], nodes[245],  nodes[1536]);
    nmos (nodes[558], nodes[985],  nodes[1536]);
    nmos (nodes[682], nodes[558],  nodes[1536]);
    nmos (nodes[665], nodes[558],  nodes[1536]);
    nmos (nodes[271], nodes[558],  nodes[1536]);
    nmos (nodes[552], nodes[558],  nodes[1536]);
    nmos (nodes[558], nodes[1623],  nodes[1536]);
    nmos (nodes[558], nodes[403],  nodes[1536]);
    nmos (nodes[558], nodes[1273],  nodes[1536]);
    nmos (nodes[1337], nodes[558],  nodes[1536]);
    nmos (nodes[1355], nodes[558],  nodes[1536]);
    nmos (nodes[787], nodes[558],  nodes[1536]);
    nmos (nodes[575], nodes[558],  nodes[1536]);
    nmos (nodes[257], nodes[558],  nodes[1536]);
    nmos (nodes[558], nodes[179],  nodes[1536]);
    nmos (nodes[558], nodes[131],  nodes[1536]);
    nmos (nodes[558], nodes[1420],  nodes[1536]);
    nmos (nodes[1342], nodes[558],  nodes[1536]);
    nmos (nodes[4], nodes[558],  nodes[1536]);
    nmos (nodes[1396], nodes[558],  nodes[1536]);
    nmos (nodes[167], nodes[558],  nodes[1536]);
    nmos (nodes[303], nodes[558],  nodes[1536]);
    nmos (nodes[558], nodes[1504],  nodes[1536]);
    nmos (nodes[558], nodes[1721],  nodes[1536]);
    nmos (nodes[558], nodes[1074],  nodes[1536]);
    nmos (nodes[1478], nodes[558],  nodes[1536]);
    nmos (nodes[594], nodes[558],  nodes[1536]);
    nmos (nodes[1292], nodes[558],  nodes[1536]);
    nmos (nodes[1114], nodes[558],  nodes[1536]);
    nmos (nodes[1476], nodes[558],  nodes[1536]);
    nmos (nodes[558], nodes[1226],  nodes[1536]);
    nmos (nodes[558], nodes[1419],  nodes[1536]);
    nmos (nodes[1491], nodes[573],  nodes[943]);
    nmos (nodes[272], nodes[558],  nodes[236]);
    nmos (nodes[299], nodes[558],  nodes[587]);
    nmos (nodes[558], nodes[1466],  nodes[337]);
    nmos (nodes[558], nodes[1601],  nodes[337]);
    nmos (nodes[1173], nodes[558],  nodes[337]);
    nmos (nodes[1562], nodes[558],  nodes[337]);
    nmos (nodes[1543], nodes[558],  nodes[337]);
    nmos (nodes[1540], nodes[558],  nodes[337]);
    nmos (nodes[245], nodes[558],  nodes[337]);
    nmos (nodes[558], nodes[985],  nodes[337]);
    nmos (nodes[558], nodes[682],  nodes[337]);
    nmos (nodes[558], nodes[665],  nodes[337]);
    nmos (nodes[286], nodes[558],  nodes[337]);
    nmos (nodes[271], nodes[558],  nodes[337]);
    nmos (nodes[370], nodes[558],  nodes[337]);
    nmos (nodes[403], nodes[558],  nodes[337]);
    nmos (nodes[804], nodes[558],  nodes[337]);
    nmos (nodes[558], nodes[712],  nodes[337]);
    nmos (nodes[558], nodes[546],  nodes[337]);
    nmos (nodes[558], nodes[776],  nodes[337]);
    nmos (nodes[257], nodes[558],  nodes[337]);
    nmos (nodes[179], nodes[558],  nodes[337]);
    nmos (nodes[1420], nodes[558],  nodes[337]);
    nmos (nodes[4], nodes[558],  nodes[337]);
    nmos (nodes[558], nodes[167],  nodes[337]);
    nmos (nodes[558], nodes[303],  nodes[337]);
    nmos (nodes[558], nodes[1504],  nodes[337]);
    nmos (nodes[558], nodes[487],  nodes[337]);
    nmos (nodes[579], nodes[558],  nodes[337]);
    nmos (nodes[145], nodes[558],  nodes[337]);
    nmos (nodes[259], nodes[558],  nodes[337]);
    nmos (nodes[517], nodes[558],  nodes[337]);
    nmos (nodes[558], nodes[352],  nodes[337]);
    nmos (nodes[558], nodes[750],  nodes[337]);
    nmos (nodes[558], nodes[528],  nodes[337]);
    nmos (nodes[558], nodes[691],  nodes[337]);
    nmos (nodes[1646], nodes[558],  nodes[337]);
    nmos (nodes[1114], nodes[558],  nodes[337]);
    nmos (nodes[1476], nodes[558],  nodes[337]);
    nmos (nodes[1226], nodes[558],  nodes[337]);
    nmos (nodes[558], nodes[1665],  nodes[337]);
    nmos (nodes[558], nodes[840],  nodes[337]);
    nmos (nodes[558], nodes[1164],  nodes[337]);
    nmos (nodes[848], nodes[473],  nodes[943]);
    nmos (nodes[389], nodes[614],  nodes[943]);
    nmos (nodes[249], nodes[558],  nodes[1359]);
    nmos (nodes[1081], nodes[960],  nodes[943]);
    nmos (nodes[558], nodes[1154],  nodes[248]);
    nmos (nodes[558], nodes[180],  nodes[248]);
    nmos (nodes[1367], nodes[558],  nodes[1202]);
    nmos (nodes[57], nodes[558],  nodes[1202]);
    nmos (nodes[620], nodes[558],  nodes[307]);
    nmos (nodes[256], nodes[558],  nodes[784]);
    nmos (nodes[278], nodes[558],  nodes[1551]);
    nmos (nodes[558], nodes[171],  nodes[567]);
    nmos (nodes[558], nodes[1026],  nodes[567]);
    nmos (nodes[322], nodes[657],  nodes[567]);
    nmos (nodes[8], nodes[558],  nodes[551]);
    nmos (nodes[1125], nodes[1620],  nodes[943]);
    nmos (nodes[558], nodes[1297],  nodes[558]);
    nmos (nodes[558], nodes[1275],  nodes[832]);
    nmos (nodes[558], nodes[437],  nodes[491]);
    nmos (nodes[558], nodes[642],  nodes[1502]);
    nmos (nodes[558], nodes[951],  nodes[1502]);
    nmos (nodes[657], nodes[1152],  nodes[1502]);
    nmos (nodes[558], nodes[744],  nodes[892]);
    nmos (nodes[696], nodes[911],  nodes[79]);
    nmos (nodes[893], nodes[277],  nodes[943]);
    nmos (nodes[558], nodes[1257],  nodes[412]);
    nmos (nodes[262], nodes[1189],  nodes[1714]);
    nmos (nodes[558], nodes[177],  nodes[1241]);
    nmos (nodes[351], nodes[558],  nodes[833]);
    nmos (nodes[1541], nodes[558],  nodes[43]);
    nmos (nodes[91], nodes[558],  nodes[1529]);
    nmos (nodes[11], nodes[558],  nodes[167]);
    nmos (nodes[1395], nodes[854],  nodes[710]);
    nmos (nodes[558], nodes[1290],  nodes[1126]);
    nmos (nodes[986], nodes[1556],  nodes[699]);
    nmos (nodes[558], nodes[867],  nodes[699]);
    nmos (nodes[558], nodes[1649],  nodes[1057]);
    nmos (nodes[1538], nodes[558],  nodes[1070]);
    nmos (nodes[558], nodes[1334],  nodes[1070]);
    nmos (nodes[200], nodes[558],  nodes[1070]);
    nmos (nodes[558], nodes[382],  nodes[1112]);
    nmos (nodes[558], nodes[1233],  nodes[1112]);
    nmos (nodes[558], nodes[84],  nodes[1112]);
    nmos (nodes[558], nodes[1543],  nodes[1112]);
    nmos (nodes[558], nodes[76],  nodes[1112]);
    nmos (nodes[558], nodes[1658],  nodes[1112]);
    nmos (nodes[558], nodes[786],  nodes[1112]);
    nmos (nodes[558], nodes[1664],  nodes[1112]);
    nmos (nodes[558], nodes[1482],  nodes[1112]);
    nmos (nodes[558], nodes[286],  nodes[1112]);
    nmos (nodes[558], nodes[271],  nodes[1112]);
    nmos (nodes[558], nodes[370],  nodes[1112]);
    nmos (nodes[558], nodes[552],  nodes[1112]);
    nmos (nodes[558], nodes[1612],  nodes[1112]);
    nmos (nodes[558], nodes[1487],  nodes[1112]);
    nmos (nodes[558], nodes[784],  nodes[1112]);
    nmos (nodes[558], nodes[764],  nodes[1112]);
    nmos (nodes[558], nodes[1057],  nodes[1112]);
    nmos (nodes[558], nodes[1582],  nodes[1112]);
    nmos (nodes[558], nodes[1031],  nodes[1112]);
    nmos (nodes[558], nodes[804],  nodes[1112]);
    nmos (nodes[558], nodes[1311],  nodes[1112]);
    nmos (nodes[558], nodes[1428],  nodes[1112]);
    nmos (nodes[558], nodes[1520],  nodes[1112]);
    nmos (nodes[558], nodes[1259],  nodes[1112]);
    nmos (nodes[558], nodes[857],  nodes[1112]);
    nmos (nodes[558], nodes[712],  nodes[1112]);
    nmos (nodes[558], nodes[1337],  nodes[1112]);
    nmos (nodes[558], nodes[1381],  nodes[1112]);
    nmos (nodes[558], nodes[776],  nodes[1112]);
    nmos (nodes[558], nodes[157],  nodes[1112]);
    nmos (nodes[558], nodes[1324],  nodes[1112]);
    nmos (nodes[558], nodes[179],  nodes[1112]);
    nmos (nodes[558], nodes[131],  nodes[1112]);
    nmos (nodes[558], nodes[4],  nodes[1112]);
    nmos (nodes[558], nodes[1396],  nodes[1112]);
    nmos (nodes[558], nodes[167],  nodes[1112]);
    nmos (nodes[558], nodes[303],  nodes[1112]);
    nmos (nodes[558], nodes[1086],  nodes[1112]);
    nmos (nodes[558], nodes[1074],  nodes[1112]);
    nmos (nodes[558], nodes[487],  nodes[1112]);
    nmos (nodes[558], nodes[579],  nodes[1112]);
    nmos (nodes[558], nodes[0],  nodes[1112]);
    nmos (nodes[558], nodes[1478],  nodes[1112]);
    nmos (nodes[558], nodes[594],  nodes[1112]);
    nmos (nodes[558], nodes[1210],  nodes[1112]);
    nmos (nodes[558], nodes[1557],  nodes[1112]);
    nmos (nodes[558], nodes[259],  nodes[1112]);
    nmos (nodes[558], nodes[1052],  nodes[1112]);
    nmos (nodes[558], nodes[791],  nodes[1112]);
    nmos (nodes[558], nodes[352],  nodes[1112]);
    nmos (nodes[558], nodes[750],  nodes[1112]);
    nmos (nodes[558], nodes[932],  nodes[1112]);
    nmos (nodes[558], nodes[1589],  nodes[1112]);
    nmos (nodes[558], nodes[446],  nodes[1112]);
    nmos (nodes[558], nodes[528],  nodes[1112]);
    nmos (nodes[558], nodes[309],  nodes[1112]);
    nmos (nodes[558], nodes[1430],  nodes[1112]);
    nmos (nodes[558], nodes[1646],  nodes[1112]);
    nmos (nodes[558], nodes[1476],  nodes[1112]);
    nmos (nodes[558], nodes[1226],  nodes[1112]);
    nmos (nodes[558], nodes[1569],  nodes[1112]);
    nmos (nodes[558], nodes[950],  nodes[1112]);
    nmos (nodes[558], nodes[1665],  nodes[1112]);
    nmos (nodes[558], nodes[1710],  nodes[1112]);
    nmos (nodes[558], nodes[1050],  nodes[1112]);
    nmos (nodes[558], nodes[607],  nodes[1112]);
    nmos (nodes[558], nodes[219],  nodes[1112]);
    nmos (nodes[558], nodes[1384],  nodes[1300]);
    nmos (nodes[1016], nodes[416],  nodes[710]);
    nmos (nodes[1637], nodes[558],  nodes[276]);
    nmos (nodes[1330], nodes[586],  nodes[1544]);
    nmos (nodes[1330], nodes[586],  nodes[1544]);
    nmos (nodes[318], nodes[1607],  nodes[943]);
    nmos (nodes[1466], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[271],  nodes[1328]);
    nmos (nodes[558], nodes[370],  nodes[1328]);
    nmos (nodes[552], nodes[558],  nodes[1328]);
    nmos (nodes[1612], nodes[558],  nodes[1328]);
    nmos (nodes[1487], nodes[558],  nodes[1328]);
    nmos (nodes[784], nodes[558],  nodes[1328]);
    nmos (nodes[244], nodes[558],  nodes[1328]);
    nmos (nodes[1623], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[764],  nodes[1328]);
    nmos (nodes[558], nodes[403],  nodes[1328]);
    nmos (nodes[1582], nodes[558],  nodes[1328]);
    nmos (nodes[1031], nodes[558],  nodes[1328]);
    nmos (nodes[804], nodes[558],  nodes[1328]);
    nmos (nodes[1311], nodes[558],  nodes[1328]);
    nmos (nodes[1520], nodes[558],  nodes[1328]);
    nmos (nodes[857], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[712],  nodes[1328]);
    nmos (nodes[1381], nodes[558],  nodes[1328]);
    nmos (nodes[546], nodes[558],  nodes[1328]);
    nmos (nodes[776], nodes[558],  nodes[1328]);
    nmos (nodes[157], nodes[558],  nodes[1328]);
    nmos (nodes[1243], nodes[558],  nodes[1328]);
    nmos (nodes[1324], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[131],  nodes[1328]);
    nmos (nodes[558], nodes[1396],  nodes[1328]);
    nmos (nodes[303], nodes[558],  nodes[1328]);
    nmos (nodes[1504], nodes[558],  nodes[1328]);
    nmos (nodes[1086], nodes[558],  nodes[1328]);
    nmos (nodes[1074], nodes[558],  nodes[1328]);
    nmos (nodes[1246], nodes[558],  nodes[1328]);
    nmos (nodes[487], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[579],  nodes[1328]);
    nmos (nodes[558], nodes[0],  nodes[1328]);
    nmos (nodes[1478], nodes[558],  nodes[1328]);
    nmos (nodes[594], nodes[558],  nodes[1328]);
    nmos (nodes[1557], nodes[558],  nodes[1328]);
    nmos (nodes[259], nodes[558],  nodes[1328]);
    nmos (nodes[1052], nodes[558],  nodes[1328]);
    nmos (nodes[791], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[352],  nodes[1328]);
    nmos (nodes[558], nodes[750],  nodes[1328]);
    nmos (nodes[932], nodes[558],  nodes[1328]);
    nmos (nodes[1589], nodes[558],  nodes[1328]);
    nmos (nodes[446], nodes[558],  nodes[1328]);
    nmos (nodes[528], nodes[558],  nodes[1328]);
    nmos (nodes[309], nodes[558],  nodes[1328]);
    nmos (nodes[1430], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[691],  nodes[1328]);
    nmos (nodes[558], nodes[1292],  nodes[1328]);
    nmos (nodes[1646], nodes[558],  nodes[1328]);
    nmos (nodes[1114], nodes[558],  nodes[1328]);
    nmos (nodes[1476], nodes[558],  nodes[1328]);
    nmos (nodes[1226], nodes[558],  nodes[1328]);
    nmos (nodes[1569], nodes[558],  nodes[1328]);
    nmos (nodes[1665], nodes[558],  nodes[1328]);
    nmos (nodes[558], nodes[1050],  nodes[1328]);
    nmos (nodes[1174], nodes[558],  nodes[1328]);
    nmos (nodes[1310], nodes[558],  nodes[1063]);
    nmos (nodes[657], nodes[672],  nodes[963]);
    nmos (nodes[846], nodes[558],  nodes[840]);
    nmos (nodes[187], nodes[558],  nodes[1131]);
    nmos (nodes[802], nodes[566],  nodes[243]);
    nmos (nodes[558], nodes[516],  nodes[216]);
    nmos (nodes[558], nodes[1610],  nodes[216]);
    nmos (nodes[1046], nodes[558],  nodes[1299]);
    nmos (nodes[558], nodes[389],  nodes[1107]);
    nmos (nodes[107], nodes[416],  nodes[639]);
    nmos (nodes[1334], nodes[558],  nodes[1007]);
    nmos (nodes[754], nodes[558],  nodes[1673]);
    nmos (nodes[707], nodes[1636],  nodes[639]);
    nmos (nodes[558], nodes[1484],  nodes[573]);
    nmos (nodes[1013], nodes[558],  nodes[1241]);
    nmos (nodes[1217], nodes[558],  nodes[1241]);
    nmos (nodes[1157], nodes[558],  nodes[291]);
    nmos (nodes[1564], nodes[657],  nodes[291]);
    nmos (nodes[558], nodes[1225],  nodes[1524]);
    nmos (nodes[10], nodes[558],  nodes[1721]);
    nmos (nodes[1488], nodes[558],  nodes[278]);
    nmos (nodes[1278], nodes[558],  nodes[462]);
    nmos (nodes[558], nodes[725],  nodes[599]);
    nmos (nodes[558], nodes[441],  nodes[692]);
    nmos (nodes[657], nodes[325],  nodes[692]);
    nmos (nodes[300], nodes[558],  nodes[1259]);
    nmos (nodes[558], nodes[1350],  nodes[760]);
    nmos (nodes[458], nodes[558],  nodes[1473]);
    nmos (nodes[558], nodes[27],  nodes[820]);
    nmos (nodes[558], nodes[917],  nodes[383]);
    nmos (nodes[386], nodes[558],  nodes[622]);
    nmos (nodes[558], nodes[1649],  nodes[248]);
    nmos (nodes[1366], nodes[472],  nodes[16]);
    nmos (nodes[850], nodes[558],  nodes[899]);
    nmos (nodes[147], nodes[558],  nodes[353]);
    nmos (nodes[147], nodes[558],  nodes[353]);
    nmos (nodes[347], nodes[558],  nodes[1385]);
    nmos (nodes[1087], nodes[1132],  nodes[710]);
    nmos (nodes[558], nodes[1180],  nodes[248]);
    nmos (nodes[188], nodes[1373],  nodes[943]);
    nmos (nodes[558], nodes[486],  nodes[817]);
    nmos (nodes[963], nodes[657],  nodes[997]);
    nmos (nodes[558], nodes[1523],  nodes[997]);
    nmos (nodes[558], nodes[635],  nodes[997]);
    nmos (nodes[558], nodes[859],  nodes[225]);
    nmos (nodes[558], nodes[136],  nodes[640]);
    nmos (nodes[558], nodes[860],  nodes[640]);
    nmos (nodes[558], nodes[1021],  nodes[155]);
    nmos (nodes[558], nodes[425],  nodes[155]);
    nmos (nodes[1555], nodes[558],  nodes[440]);
    nmos (nodes[558], nodes[1686],  nodes[432]);
    nmos (nodes[558], nodes[1097],  nodes[432]);
    nmos (nodes[672], nodes[558],  nodes[635]);
    nmos (nodes[558], nodes[672],  nodes[635]);
    nmos (nodes[672], nodes[558],  nodes[635]);
    nmos (nodes[558], nodes[672],  nodes[635]);
    nmos (nodes[672], nodes[558],  nodes[635]);
    nmos (nodes[558], nodes[672],  nodes[635]);
    nmos (nodes[558], nodes[672],  nodes[635]);
    nmos (nodes[1534], nodes[558],  nodes[43]);
    nmos (nodes[558], nodes[1330],  nodes[967]);
    nmos (nodes[558], nodes[721],  nodes[181]);
    nmos (nodes[683], nodes[1225],  nodes[943]);
    nmos (nodes[630], nodes[558],  nodes[726]);
    nmos (nodes[1191], nodes[558],  nodes[1195]);
    nmos (nodes[657], nodes[1254],  nodes[1195]);
    nmos (nodes[558], nodes[1055],  nodes[771]);
    nmos (nodes[558], nodes[251],  nodes[221]);
    nmos (nodes[251], nodes[558],  nodes[221]);
    nmos (nodes[372], nodes[558],  nodes[248]);
    nmos (nodes[1085], nodes[1365],  nodes[248]);
    nmos (nodes[92], nodes[359],  nodes[943]);
    nmos (nodes[756], nodes[626],  nodes[710]);
    nmos (nodes[823], nodes[457],  nodes[710]);
    nmos (nodes[741], nodes[558],  nodes[255]);
    nmos (nodes[657], nodes[148],  nodes[1140]);
    nmos (nodes[558], nodes[1634],  nodes[1288]);
    nmos (nodes[1040], nodes[558],  nodes[383]);
    nmos (nodes[558], nodes[1040],  nodes[383]);
    nmos (nodes[699], nodes[558],  nodes[1637]);
    nmos (nodes[1495], nodes[1445],  nodes[270]);
    nmos (nodes[1552], nodes[558],  nodes[1593]);
    nmos (nodes[657], nodes[362],  nodes[1593]);
    nmos (nodes[957], nodes[1525],  nodes[1666]);
    nmos (nodes[953], nodes[250],  nodes[1666]);
    nmos (nodes[740], nodes[701],  nodes[1666]);
    nmos (nodes[1071], nodes[884],  nodes[1666]);
    nmos (nodes[296], nodes[308],  nodes[1666]);
    nmos (nodes[277], nodes[1469],  nodes[1666]);
    nmos (nodes[722], nodes[1459],  nodes[1666]);
    nmos (nodes[177], nodes[304],  nodes[1666]);
    nmos (nodes[256], nodes[558],  nodes[341]);
    nmos (nodes[428], nodes[1558],  nodes[16]);
    nmos (nodes[591], nodes[252],  nodes[691]);
    nmos (nodes[1672], nodes[558],  nodes[558]);
    nmos (nodes[558], nodes[1053],  nodes[439]);
    nmos (nodes[786], nodes[558],  nodes[156]);
    nmos (nodes[1664], nodes[558],  nodes[156]);
    nmos (nodes[1482], nodes[558],  nodes[156]);
    nmos (nodes[1243], nodes[558],  nodes[156]);
    nmos (nodes[822], nodes[558],  nodes[156]);
    nmos (nodes[558], nodes[1324],  nodes[156]);
    nmos (nodes[1646], nodes[558],  nodes[156]);
    nmos (nodes[558], nodes[1155],  nodes[156]);
    nmos (nodes[301], nodes[558],  nodes[156]);
    nmos (nodes[950], nodes[558],  nodes[156]);
    nmos (nodes[1665], nodes[558],  nodes[156]);
    nmos (nodes[1710], nodes[558],  nodes[156]);
    nmos (nodes[657], nodes[1302],  nodes[943]);
    nmos (nodes[1], nodes[1694],  nodes[943]);
    nmos (nodes[1403], nodes[54],  nodes[874]);
    nmos (nodes[137], nodes[558],  nodes[1120]);
    nmos (nodes[558], nodes[1171],  nodes[558]);
    nmos (nodes[558], nodes[744],  nodes[833]);
    nmos (nodes[558], nodes[218],  nodes[368]);
    nmos (nodes[1707], nodes[319],  nodes[623]);
    nmos (nodes[558], nodes[388],  nodes[623]);
    nmos (nodes[558], nodes[1368],  nodes[1578]);
    nmos (nodes[476], nodes[558],  nodes[1027]);
    nmos (nodes[558], nodes[368],  nodes[1589]);
    nmos (nodes[558], nodes[104],  nodes[1589]);
    nmos (nodes[1096], nodes[558],  nodes[153]);
    nmos (nodes[558], nodes[1352],  nodes[440]);
    nmos (nodes[558], nodes[104],  nodes[440]);
    nmos (nodes[558], nodes[812],  nodes[440]);
    nmos (nodes[962], nodes[558],  nodes[1585]);
    nmos (nodes[558], nodes[1489],  nodes[1398]);
    nmos (nodes[1106], nodes[1103],  nodes[258]);
    nmos (nodes[558], nodes[1347],  nodes[979]);
    nmos (nodes[1464], nodes[558],  nodes[370]);
    nmos (nodes[1671], nodes[558],  nodes[955]);
    nmos (nodes[558], nodes[911],  nodes[1343]);
    nmos (nodes[434], nodes[558],  nodes[790]);
    nmos (nodes[70], nodes[558],  nodes[1054]);
    nmos (nodes[1106], nodes[558],  nodes[1543]);
    nmos (nodes[558], nodes[320],  nodes[1150]);
    nmos (nodes[488], nodes[1108],  nodes[283]);
    nmos (nodes[1608], nodes[657],  nodes[775]);
    nmos (nodes[558], nodes[1423],  nodes[775]);
    nmos (nodes[558], nodes[869],  nodes[775]);
    nmos (nodes[481], nodes[1473],  nodes[283]);
    nmos (nodes[558], nodes[340],  nodes[1164]);
    nmos (nodes[1382], nodes[558],  nodes[248]);
    nmos (nodes[1053], nodes[673],  nodes[575]);
    nmos (nodes[927], nodes[703],  nodes[879]);
    nmos (nodes[558], nodes[931],  nodes[415]);
    nmos (nodes[558], nodes[1375],  nodes[88]);
    nmos (nodes[558], nodes[771],  nodes[1110]);
    nmos (nodes[1388], nodes[965],  nodes[1506]);
    nmos (nodes[558], nodes[295],  nodes[1506]);
    nmos (nodes[7], nodes[558],  nodes[353]);
    nmos (nodes[7], nodes[558],  nodes[353]);
    nmos (nodes[466], nodes[558],  nodes[353]);
    nmos (nodes[558], nodes[920],  nodes[73]);
    nmos (nodes[558], nodes[651],  nodes[65]);
    nmos (nodes[902], nodes[248],  nodes[710]);
    nmos (nodes[558], nodes[1182],  nodes[1384]);
    nmos (nodes[895], nodes[1675],  nodes[943]);
    nmos (nodes[558], nodes[674],  nodes[25]);
    nmos (nodes[829], nodes[1588],  nodes[943]);
    nmos (nodes[1281], nodes[894],  nodes[943]);
    nmos (nodes[1075], nodes[369],  nodes[943]);
    nmos (nodes[1234], nodes[929],  nodes[943]);
    nmos (nodes[1223], nodes[558],  nodes[688]);
    nmos (nodes[1537], nodes[1638],  nodes[943]);
    nmos (nodes[716], nodes[701],  nodes[110]);
    nmos (nodes[558], nodes[1716],  nodes[510]);
    nmos (nodes[558], nodes[161],  nodes[1113]);
    nmos (nodes[558], nodes[1382],  nodes[861]);
    nmos (nodes[1068], nodes[558],  nodes[1247]);
    nmos (nodes[1591], nodes[1591],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[1591], nodes[558],  nodes[471]);
    nmos (nodes[558], nodes[1591],  nodes[471]);
    nmos (nodes[1325], nodes[558],  nodes[353]);
    nmos (nodes[1325], nodes[558],  nodes[353]);
    nmos (nodes[769], nodes[558],  nodes[353]);
    nmos (nodes[657], nodes[1467],  nodes[358]);
    nmos (nodes[1094], nodes[463],  nodes[710]);
    nmos (nodes[1620], nodes[1590],  nodes[879]);
    nmos (nodes[1368], nodes[558],  nodes[645]);
    nmos (nodes[1275], nodes[558],  nodes[248]);
    nmos (nodes[1267], nodes[558],  nodes[52]);
    nmos (nodes[514], nodes[494],  nodes[710]);
    nmos (nodes[558], nodes[279],  nodes[954]);
    nmos (nodes[558], nodes[367],  nodes[954]);
    nmos (nodes[1427], nodes[558],  nodes[236]);
    nmos (nodes[1464], nodes[558],  nodes[271]);
    nmos (nodes[1496], nodes[558],  nodes[114]);
    nmos (nodes[843], nodes[1251],  nodes[943]);
    nmos (nodes[1519], nodes[558],  nodes[1437]);
    nmos (nodes[1447], nodes[262],  nodes[710]);
    nmos (nodes[1196], nodes[558],  nodes[522]);
    nmos (nodes[153], nodes[246],  nodes[639]);
    nmos (nodes[790], nodes[558],  nodes[691]);
    nmos (nodes[558], nodes[1601],  nodes[1182]);
    nmos (nodes[558], nodes[258],  nodes[1182]);
    nmos (nodes[558], nodes[665],  nodes[1182]);
    nmos (nodes[558], nodes[764],  nodes[1182]);
    nmos (nodes[558], nodes[1057],  nodes[1182]);
    nmos (nodes[558], nodes[1381],  nodes[1182]);
    nmos (nodes[558], nodes[303],  nodes[1182]);
    nmos (nodes[558], nodes[285],  nodes[1182]);
    nmos (nodes[558], nodes[594],  nodes[1182]);
    nmos (nodes[558], nodes[1052],  nodes[1182]);
    nmos (nodes[558], nodes[1589],  nodes[1182]);
    nmos (nodes[558], nodes[309],  nodes[1182]);
    nmos (nodes[558], nodes[1646],  nodes[1182]);
    nmos (nodes[558], nodes[904],  nodes[1182]);
    nmos (nodes[558], nodes[1476],  nodes[1182]);
    nmos (nodes[558], nodes[950],  nodes[1182]);
    nmos (nodes[607], nodes[558],  nodes[1182]);
    nmos (nodes[558], nodes[219],  nodes[1182]);
    nmos (nodes[984], nodes[558],  nodes[943]);
    nmos (nodes[549], nodes[558],  nodes[943]);
    nmos (nodes[437], nodes[558],  nodes[943]);
    nmos (nodes[859], nodes[558],  nodes[943]);
    nmos (nodes[1068], nodes[558],  nodes[943]);
    nmos (nodes[654], nodes[558],  nodes[943]);
    nmos (nodes[558], nodes[874],  nodes[943]);
    nmos (nodes[1167], nodes[558],  nodes[984]);
    nmos (nodes[792], nodes[851],  nodes[710]);
    nmos (nodes[1248], nodes[558],  nodes[984]);
    nmos (nodes[1142], nodes[558],  nodes[984]);
    nmos (nodes[1627], nodes[558],  nodes[984]);
    nmos (nodes[530], nodes[558],  nodes[984]);
    nmos (nodes[510], nodes[558],  nodes[1052]);
    nmos (nodes[134], nodes[558],  nodes[1052]);
    nmos (nodes[558], nodes[105],  nodes[1165]);
    nmos (nodes[942], nodes[558],  nodes[1165]);
    nmos (nodes[945], nodes[945],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[945], nodes[558],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[558], nodes[945],  nodes[37]);
    nmos (nodes[945], nodes[558],  nodes[37]);
    nmos (nodes[558], nodes[36],  nodes[8]);
    nmos (nodes[558], nodes[150],  nodes[8]);
    nmos (nodes[333], nodes[1030],  nodes[570]);
    nmos (nodes[558], nodes[591],  nodes[1258]);
    nmos (nodes[657], nodes[684],  nodes[943]);
    nmos (nodes[1649], nodes[558],  nodes[1259]);
    nmos (nodes[448], nodes[1724],  nodes[943]);
    nmos (nodes[1598], nodes[558],  nodes[685]);
    nmos (nodes[1060], nodes[558],  nodes[1238]);
    nmos (nodes[957], nodes[371],  nodes[921]);
    nmos (nodes[250], nodes[965],  nodes[921]);
    nmos (nodes[740], nodes[22],  nodes[921]);
    nmos (nodes[1071], nodes[274],  nodes[921]);
    nmos (nodes[296], nodes[651],  nodes[921]);
    nmos (nodes[277], nodes[486],  nodes[921]);
    nmos (nodes[1197], nodes[722],  nodes[921]);
    nmos (nodes[532], nodes[304],  nodes[921]);
    nmos (nodes[1288], nodes[1376],  nodes[710]);
    nmos (nodes[327], nodes[558],  nodes[1569]);
    nmos (nodes[558], nodes[640],  nodes[988]);
    nmos (nodes[828], nodes[34],  nodes[943]);
    nmos (nodes[1188], nodes[657],  nodes[943]);
    nmos (nodes[2], nodes[558],  nodes[151]);
    nmos (nodes[558], nodes[72],  nodes[1326]);
    nmos (nodes[597], nodes[1339],  nodes[710]);
    nmos (nodes[834], nodes[558],  nodes[402]);
    nmos (nodes[558], nodes[436],  nodes[485]);
    nmos (nodes[558], nodes[809],  nodes[361]);
    nmos (nodes[509], nodes[442],  nodes[943]);
    nmos (nodes[564], nodes[558],  nodes[1025]);
    nmos (nodes[1601], nodes[558],  nodes[1320]);
    nmos (nodes[382], nodes[558],  nodes[1320]);
    nmos (nodes[1173], nodes[558],  nodes[1320]);
    nmos (nodes[1233], nodes[558],  nodes[1320]);
    nmos (nodes[558], nodes[1562],  nodes[1320]);
    nmos (nodes[1543], nodes[558],  nodes[1320]);
    nmos (nodes[76], nodes[558],  nodes[1320]);
    nmos (nodes[1658], nodes[558],  nodes[1320]);
    nmos (nodes[1540], nodes[558],  nodes[1320]);
    nmos (nodes[245], nodes[558],  nodes[1320]);
    nmos (nodes[985], nodes[558],  nodes[1320]);
    nmos (nodes[786], nodes[558],  nodes[1320]);
    nmos (nodes[558], nodes[1664],  nodes[1320]);
    nmos (nodes[682], nodes[558],  nodes[1320]);
    nmos (nodes[1482], nodes[558],  nodes[1320]);
    nmos (nodes[665], nodes[558],  nodes[1320]);
    nmos (nodes[286], nodes[558],  nodes[1320]);
    nmos (nodes[324], nodes[558],  nodes[1320]);
    nmos (nodes[1337], nodes[558],  nodes[1320]);
    nmos (nodes[1355], nodes[558],  nodes[1320]);
    nmos (nodes[787], nodes[558],  nodes[1320]);
    nmos (nodes[257], nodes[558],  nodes[1320]);
    nmos (nodes[179], nodes[558],  nodes[1320]);
    nmos (nodes[1420], nodes[558],  nodes[1320]);
    nmos (nodes[4], nodes[558],  nodes[1320]);
    nmos (nodes[167], nodes[558],  nodes[1320]);
    nmos (nodes[145], nodes[558],  nodes[1320]);
    nmos (nodes[517], nodes[558],  nodes[1320]);
    nmos (nodes[301], nodes[558],  nodes[1320]);
    nmos (nodes[950], nodes[558],  nodes[1320]);
    nmos (nodes[558], nodes[1710],  nodes[1320]);
    nmos (nodes[558], nodes[1419],  nodes[1320]);
    nmos (nodes[1164], nodes[558],  nodes[1320]);
    nmos (nodes[624], nodes[977],  nodes[1068]);
    nmos (nodes[79], nodes[558],  nodes[236]);
    nmos (nodes[558], nodes[1003],  nodes[1023]);
    nmos (nodes[924], nodes[1425],  nodes[1023]);
    nmos (nodes[478], nodes[1645],  nodes[1068]);
    nmos (nodes[458], nodes[704],  nodes[1068]);
    nmos (nodes[558], nodes[753],  nodes[811]);
    nmos (nodes[558], nodes[753],  nodes[811]);
    nmos (nodes[127], nodes[558],  nodes[519]);
    nmos (nodes[657], nodes[135],  nodes[519]);
    nmos (nodes[558], nodes[1575],  nodes[1360]);
    nmos (nodes[252], nodes[558],  nodes[1155]);
    nmos (nodes[558], nodes[1348],  nodes[1628]);
    nmos (nodes[468], nodes[1703],  nodes[16]);
    nmos (nodes[558], nodes[366],  nodes[1074]);
    nmos (nodes[1583], nodes[308],  nodes[1063]);
    nmos (nodes[234], nodes[558],  nodes[1513]);
    nmos (nodes[384], nodes[558],  nodes[946]);
    nmos (nodes[128], nodes[558],  nodes[1653]);
    nmos (nodes[558], nodes[275],  nodes[773]);
    nmos (nodes[558], nodes[66],  nodes[376]);
    nmos (nodes[842], nodes[558],  nodes[376]);
    nmos (nodes[657], nodes[1479],  nodes[376]);
    nmos (nodes[1709], nodes[98],  nodes[943]);
    nmos (nodes[1282], nodes[558],  nodes[686]);
    nmos (nodes[645], nodes[562],  nodes[710]);
    nmos (nodes[558], nodes[1705],  nodes[467]);
    nmos (nodes[346], nodes[297],  nodes[1392]);
    nmos (nodes[284], nodes[558],  nodes[1392]);
    nmos (nodes[1227], nodes[558],  nodes[526]);
    nmos (nodes[1464], nodes[558],  nodes[552]);
    nmos (nodes[78], nodes[558],  nodes[1425]);
    nmos (nodes[142], nodes[1310],  nodes[1425]);
    nmos (nodes[1617], nodes[558],  nodes[117]);
    nmos (nodes[558], nodes[422],  nodes[92]);
    nmos (nodes[744], nodes[558],  nodes[991]);
    nmos (nodes[558], nodes[851],  nodes[1294]);
    nmos (nodes[944], nodes[197],  nodes[943]);
    nmos (nodes[1106], nodes[558],  nodes[1658]);
    nmos (nodes[1418], nodes[1684],  nodes[710]);
    nmos (nodes[558], nodes[388],  nodes[516]);
    nmos (nodes[558], nodes[1566],  nodes[1221]);
    nmos (nodes[1044], nodes[558],  nodes[812]);
    nmos (nodes[1131], nodes[1352],  nodes[943]);
    nmos (nodes[1560], nodes[558],  nodes[1355]);
    nmos (nodes[95], nodes[1375],  nodes[710]);
    nmos (nodes[1529], nodes[1089],  nodes[710]);
    nmos (nodes[946], nodes[454],  nodes[844]);
    nmos (nodes[1336], nodes[331],  nodes[129]);
    nmos (nodes[166], nodes[314],  nodes[129]);
    nmos (nodes[606], nodes[1405],  nodes[129]);
    nmos (nodes[1188], nodes[1414],  nodes[129]);
    nmos (nodes[558], nodes[1391],  nodes[352]);
    nmos (nodes[558], nodes[1352],  nodes[352]);
    nmos (nodes[1657], nodes[820],  nodes[943]);
    nmos (nodes[845], nodes[511],  nodes[553]);
    nmos (nodes[608], nodes[558],  nodes[1272]);
    nmos (nodes[123], nodes[558],  nodes[413]);
    nmos (nodes[185], nodes[558],  nodes[1142]);
    nmos (nodes[404], nodes[558],  nodes[1142]);
    nmos (nodes[558], nodes[21],  nodes[43]);
    nmos (nodes[944], nodes[558],  nodes[1449]);
    nmos (nodes[558], nodes[337],  nodes[1675]);
    nmos (nodes[1091], nodes[363],  nodes[16]);
    nmos (nodes[1717], nodes[558],  nodes[1233]);
    nmos (nodes[558], nodes[885],  nodes[384]);
    nmos (nodes[558], nodes[550],  nodes[384]);
    nmos (nodes[598], nodes[176],  nodes[943]);
    nmos (nodes[1653], nodes[1592],  nodes[943]);
    nmos (nodes[891], nodes[558],  nodes[943]);
    nmos (nodes[1562], nodes[558],  nodes[702]);
    nmos (nodes[558], nodes[1543],  nodes[702]);
    nmos (nodes[558], nodes[76],  nodes[702]);
    nmos (nodes[558], nodes[1540],  nodes[702]);
    nmos (nodes[558], nodes[245],  nodes[702]);
    nmos (nodes[558], nodes[985],  nodes[702]);
    nmos (nodes[558], nodes[786],  nodes[702]);
    nmos (nodes[558], nodes[682],  nodes[702]);
    nmos (nodes[558], nodes[244],  nodes[702]);
    nmos (nodes[558], nodes[324],  nodes[702]);
    nmos (nodes[1466], nodes[558],  nodes[702]);
    nmos (nodes[558], nodes[546],  nodes[702]);
    nmos (nodes[558], nodes[1324],  nodes[702]);
    nmos (nodes[558], nodes[179],  nodes[702]);
    nmos (nodes[558], nodes[1396],  nodes[702]);
    nmos (nodes[558], nodes[167],  nodes[702]);
    nmos (nodes[558], nodes[1074],  nodes[702]);
    nmos (nodes[558], nodes[1246],  nodes[702]);
    nmos (nodes[558], nodes[53],  nodes[702]);
    nmos (nodes[558], nodes[691],  nodes[702]);
    nmos (nodes[558], nodes[1665],  nodes[702]);
    nmos (nodes[191], nodes[558],  nodes[248]);
    nmos (nodes[1275], nodes[558],  nodes[778]);
    nmos (nodes[558], nodes[687],  nodes[31]);
    nmos (nodes[42], nodes[657],  nodes[444]);
    nmos (nodes[558], nodes[1196],  nodes[1228]);
    nmos (nodes[657], nodes[148],  nodes[1140]);
    nmos (nodes[1036], nodes[67],  nodes[943]);
    nmos (nodes[558], nodes[1236],  nodes[1632]);
    nmos (nodes[558], nodes[1220],  nodes[1632]);
    nmos (nodes[558], nodes[1498],  nodes[163]);
    nmos (nodes[558], nodes[903],  nodes[163]);
    nmos (nodes[558], nodes[1576],  nodes[1620]);
    nmos (nodes[862], nodes[1011],  nodes[943]);
    nmos (nodes[222], nodes[1687],  nodes[710]);
    nmos (nodes[1625], nodes[299],  nodes[710]);
    nmos (nodes[169], nodes[1008],  nodes[943]);
    nmos (nodes[558], nodes[1714],  nodes[1321]);
    nmos (nodes[558], nodes[1103],  nodes[1244]);
    nmos (nodes[558], nodes[620],  nodes[1433]);
    nmos (nodes[1353], nodes[254],  nodes[710]);
    nmos (nodes[1283], nodes[340],  nodes[943]);
    nmos (nodes[1023], nodes[433],  nodes[681]);
    nmos (nodes[206], nodes[430],  nodes[1446]);
    nmos (nodes[558], nodes[311],  nodes[1010]);
    nmos (nodes[558], nodes[1334],  nodes[1010]);
    nmos (nodes[534], nodes[558],  nodes[1047]);
    nmos (nodes[558], nodes[35],  nodes[796]);
    nmos (nodes[933], nodes[1407],  nodes[1262]);
    nmos (nodes[1490], nodes[296],  nodes[943]);
    nmos (nodes[928], nodes[558],  nodes[667]);
    nmos (nodes[1032], nodes[891],  nodes[284]);
    nmos (nodes[558], nodes[1070],  nodes[292]);
    nmos (nodes[558], nodes[60],  nodes[26]);
    nmos (nodes[558], nodes[1512],  nodes[26]);
    nmos (nodes[558], nodes[1173],  nodes[26]);
    nmos (nodes[558], nodes[258],  nodes[26]);
    nmos (nodes[558], nodes[245],  nodes[26]);
    nmos (nodes[558], nodes[682],  nodes[26]);
    nmos (nodes[558], nodes[492],  nodes[26]);
    nmos (nodes[558], nodes[1204],  nodes[26]);
    nmos (nodes[58], nodes[558],  nodes[26]);
    nmos (nodes[558], nodes[342],  nodes[26]);
    nmos (nodes[558], nodes[257],  nodes[26]);
    nmos (nodes[558], nodes[354],  nodes[26]);
    nmos (nodes[558], nodes[1168],  nodes[26]);
    nmos (nodes[558], nodes[1721],  nodes[26]);
    nmos (nodes[558], nodes[1239],  nodes[26]);
    nmos (nodes[461], nodes[558],  nodes[26]);
    nmos (nodes[558], nodes[447],  nodes[26]);
    nmos (nodes[558], nodes[660],  nodes[26]);
    nmos (nodes[558], nodes[1292],  nodes[26]);
    nmos (nodes[558], nodes[1114],  nodes[26]);
    nmos (nodes[558], nodes[904],  nodes[26]);
    nmos (nodes[1419], nodes[558],  nodes[26]);
    nmos (nodes[558], nodes[281],  nodes[26]);
    nmos (nodes[558], nodes[1164],  nodes[26]);
    nmos (nodes[168], nodes[558],  nodes[1651]);
    nmos (nodes[704], nodes[1242],  nodes[437]);
    nmos (nodes[1104], nodes[889],  nodes[943]);
    nmos (nodes[558], nodes[1474],  nodes[991]);
    nmos (nodes[558], nodes[48],  nodes[1247]);
    nmos (nodes[558], nodes[1331],  nodes[1247]);
    nmos (nodes[558], nodes[1039],  nodes[456]);
    nmos (nodes[558], nodes[939],  nodes[647]);
    nmos (nodes[138], nodes[825],  nodes[943]);
    nmos (nodes[558], nodes[717],  nodes[1036]);
    nmos (nodes[1650], nodes[558],  nodes[1672]);
    nmos (nodes[558], nodes[1270],  nodes[509]);
    nmos (nodes[390], nodes[558],  nodes[653]);
    nmos (nodes[1455], nodes[558],  nodes[179]);
    nmos (nodes[558], nodes[1365],  nodes[862]);
    nmos (nodes[9], nodes[657],  nodes[866]);
    nmos (nodes[558], nodes[1560],  nodes[1055]);
    nmos (nodes[558], nodes[269],  nodes[1038]);
    nmos (nodes[1019], nodes[558],  nodes[1622]);
    nmos (nodes[558], nodes[1294],  nodes[1622]);
    nmos (nodes[1491], nodes[558],  nodes[1484]);
    nmos (nodes[1374], nodes[558],  nodes[882]);
    nmos (nodes[558], nodes[306],  nodes[725]);
    nmos (nodes[558], nodes[1619],  nodes[1448]);
    nmos (nodes[858], nodes[831],  nodes[943]);
    nmos (nodes[262], nodes[1598],  nodes[1511]);
    nmos (nodes[991], nodes[1444],  nodes[1042]);
    nmos (nodes[558], nodes[1633],  nodes[172]);
    nmos (nodes[657], nodes[210],  nodes[172]);
    nmos (nodes[558], nodes[678],  nodes[1357]);
    nmos (nodes[1600], nodes[558],  nodes[1302]);
    nmos (nodes[1150], nodes[98],  nodes[1186]);
    nmos (nodes[964], nodes[558],  nodes[1533]);
    nmos (nodes[558], nodes[149],  nodes[331]);
    nmos (nodes[1522], nodes[558],  nodes[984]);
    nmos (nodes[1399], nodes[558],  nodes[1715]);
    nmos (nodes[1399], nodes[558],  nodes[1715]);
    nmos (nodes[657], nodes[1105],  nodes[1715]);
    nmos (nodes[558], nodes[726],  nodes[677]);
    nmos (nodes[558], nodes[565],  nodes[989]);
    nmos (nodes[329], nodes[558],  nodes[1022]);
    nmos (nodes[1465], nodes[558],  nodes[689]);
    nmos (nodes[796], nodes[396],  nodes[943]);
    nmos (nodes[1100], nodes[153],  nodes[943]);
    nmos (nodes[558], nodes[793],  nodes[1442]);
    nmos (nodes[109], nodes[558],  nodes[1380]);
    nmos (nodes[405], nodes[558],  nodes[967]);
    nmos (nodes[558], nodes[1312],  nodes[1693]);
    nmos (nodes[558], nodes[1604],  nodes[1601]);
    nmos (nodes[1397], nodes[558],  nodes[1601]);
    nmos (nodes[1698], nodes[558],  nodes[1247]);
    nmos (nodes[175], nodes[558],  nodes[558]);
    nmos (nodes[333], nodes[1030],  nodes[269]);
    nmos (nodes[558], nodes[1721],  nodes[603]);
    nmos (nodes[336], nodes[1483],  nodes[235]);
    nmos (nodes[1084], nodes[558],  nodes[235]);
    nmos (nodes[558], nodes[970],  nodes[149]);
    nmos (nodes[762], nodes[558],  nodes[149]);
    nmos (nodes[478], nodes[558],  nodes[892]);
    nmos (nodes[558], nodes[965],  nodes[295]);
    nmos (nodes[558], nodes[273],  nodes[791]);
    nmos (nodes[558], nodes[677],  nodes[791]);
    nmos (nodes[558], nodes[1597],  nodes[116]);
    nmos (nodes[1597], nodes[558],  nodes[116]);
    nmos (nodes[558], nodes[1597],  nodes[116]);
    nmos (nodes[966], nodes[558],  nodes[1683]);
    nmos (nodes[558], nodes[325],  nodes[441]);
    nmos (nodes[1649], nodes[558],  nodes[1109]);
    nmos (nodes[318], nodes[558],  nodes[627]);
    nmos (nodes[881], nodes[330],  nodes[538]);
    nmos (nodes[1223], nodes[558],  nodes[43]);
    nmos (nodes[558], nodes[874],  nodes[282]);
    nmos (nodes[1301], nodes[558],  nodes[33]);
    nmos (nodes[558], nodes[1517],  nodes[853]);
    nmos (nodes[558], nodes[1388],  nodes[425]);
    nmos (nodes[558], nodes[295],  nodes[425]);
    nmos (nodes[558], nodes[1584],  nodes[876]);
    nmos (nodes[833], nodes[1458],  nodes[283]);
    nmos (nodes[558], nodes[326],  nodes[1356]);
    nmos (nodes[558], nodes[637],  nodes[1318]);
    nmos (nodes[558], nodes[516],  nodes[1691]);
    nmos (nodes[401], nodes[558],  nodes[394]);
    nmos (nodes[471], nodes[558],  nodes[1415]);
    nmos (nodes[466], nodes[558],  nodes[1415]);
    nmos (nodes[698], nodes[1290],  nodes[710]);
    nmos (nodes[955], nodes[111],  nodes[943]);
    nmos (nodes[1690], nodes[62],  nodes[943]);
    nmos (nodes[1669], nodes[374],  nodes[943]);
    nmos (nodes[558], nodes[888],  nodes[675]);
    nmos (nodes[558], nodes[888],  nodes[675]);
    nmos (nodes[872], nodes[558],  nodes[697]);
    nmos (nodes[558], nodes[636],  nodes[1239]);
    nmos (nodes[106], nodes[732],  nodes[792]);
    nmos (nodes[93], nodes[558],  nodes[1005]);
    nmos (nodes[558], nodes[419],  nodes[978]);
    nmos (nodes[1320], nodes[558],  nodes[1328]);
    nmos (nodes[1688], nodes[558],  nodes[1304]);
    nmos (nodes[998], nodes[558],  nodes[828]);
    nmos (nodes[558], nodes[1145],  nodes[248]);
    nmos (nodes[558], nodes[604],  nodes[248]);
    nmos (nodes[599], nodes[533],  nodes[710]);
    nmos (nodes[694], nodes[558],  nodes[1064]);
    nmos (nodes[849], nodes[558],  nodes[321]);
    nmos (nodes[247], nodes[657],  nodes[321]);
    nmos (nodes[558], nodes[384],  nodes[1228]);
    nmos (nodes[558], nodes[384],  nodes[1228]);
    nmos (nodes[558], nodes[385],  nodes[1377]);
    nmos (nodes[1614], nodes[558],  nodes[1177]);
    nmos (nodes[300], nodes[558],  nodes[857]);
    nmos (nodes[520], nodes[558],  nodes[353]);
    nmos (nodes[520], nodes[558],  nodes[353]);
    nmos (nodes[224], nodes[558],  nodes[353]);
    nmos (nodes[558], nodes[60],  nodes[194]);
    nmos (nodes[558], nodes[1512],  nodes[194]);
    nmos (nodes[558], nodes[84],  nodes[194]);
    nmos (nodes[1623], nodes[558],  nodes[194]);
    nmos (nodes[403], nodes[558],  nodes[194]);
    nmos (nodes[1428], nodes[558],  nodes[194]);
    nmos (nodes[492], nodes[558],  nodes[194]);
    nmos (nodes[1204], nodes[558],  nodes[194]);
    nmos (nodes[558], nodes[1259],  nodes[194]);
    nmos (nodes[342], nodes[558],  nodes[194]);
    nmos (nodes[1355], nodes[558],  nodes[194]);
    nmos (nodes[787], nodes[558],  nodes[194]);
    nmos (nodes[575], nodes[558],  nodes[194]);
    nmos (nodes[558], nodes[1243],  nodes[194]);
    nmos (nodes[558], nodes[822],  nodes[194]);
    nmos (nodes[558], nodes[1420],  nodes[194]);
    nmos (nodes[1342], nodes[558],  nodes[194]);
    nmos (nodes[1504], nodes[558],  nodes[194]);
    nmos (nodes[558], nodes[1168],  nodes[194]);
    nmos (nodes[558], nodes[145],  nodes[194]);
    nmos (nodes[558], nodes[1524],  nodes[194]);
    nmos (nodes[558], nodes[1210],  nodes[194]);
    nmos (nodes[558], nodes[461],  nodes[194]);
    nmos (nodes[1155], nodes[558],  nodes[194]);
    nmos (nodes[301], nodes[558],  nodes[194]);
    nmos (nodes[1385], nodes[558],  nodes[194]);
    nmos (nodes[650], nodes[558],  nodes[558]);
    nmos (nodes[944], nodes[558],  nodes[759]);
    nmos (nodes[343], nodes[1300],  nodes[879]);
    nmos (nodes[664], nodes[558],  nodes[1006]);
    nmos (nodes[330], nodes[675],  nodes[710]);
    nmos (nodes[558], nodes[612],  nodes[353]);
    nmos (nodes[558], nodes[612],  nodes[353]);
    nmos (nodes[294], nodes[14],  nodes[943]);
    nmos (nodes[832], nodes[586],  nodes[943]);
    nmos (nodes[60], nodes[558],  nodes[1567]);
    nmos (nodes[1487], nodes[558],  nodes[1567]);
    nmos (nodes[1031], nodes[558],  nodes[1567]);
    nmos (nodes[558], nodes[1428],  nodes[1567]);
    nmos (nodes[58], nodes[558],  nodes[1567]);
    nmos (nodes[342], nodes[558],  nodes[1567]);
    nmos (nodes[558], nodes[1381],  nodes[1567]);
    nmos (nodes[579], nodes[558],  nodes[1567]);
    nmos (nodes[120], nodes[558],  nodes[1567]);
    nmos (nodes[677], nodes[558],  nodes[1567]);
    nmos (nodes[447], nodes[558],  nodes[1567]);
    nmos (nodes[660], nodes[558],  nodes[1567]);
    nmos (nodes[1430], nodes[558],  nodes[1567]);
    nmos (nodes[558], nodes[904],  nodes[1567]);
    nmos (nodes[607], nodes[558],  nodes[1567]);
    nmos (nodes[150], nodes[613],  nodes[1682]);
    nmos (nodes[1256], nodes[558],  nodes[91]);
    nmos (nodes[574], nodes[657],  nodes[91]);
    nmos (nodes[543], nodes[558],  nodes[339]);
    nmos (nodes[558], nodes[239],  nodes[595]);
    nmos (nodes[558], nodes[992],  nodes[595]);
    nmos (nodes[859], nodes[558],  nodes[1247]);
    nmos (nodes[907], nodes[676],  nodes[943]);
    nmos (nodes[1536], nodes[657],  nodes[17]);
    nmos (nodes[646], nodes[558],  nodes[17]);
    nmos (nodes[889], nodes[558],  nodes[1114]);
    nmos (nodes[558], nodes[327],  nodes[1226]);
    nmos (nodes[1661], nodes[684],  nodes[1564]);
    nmos (nodes[1095], nodes[1437],  nodes[1564]);
    nmos (nodes[87], nodes[1282],  nodes[1564]);
    nmos (nodes[1424], nodes[1242],  nodes[1564]);
    nmos (nodes[719], nodes[413],  nodes[1564]);
    nmos (nodes[558], nodes[1322],  nodes[320]);
    nmos (nodes[558], nodes[735],  nodes[320]);
    nmos (nodes[471], nodes[558],  nodes[353]);
    nmos (nodes[471], nodes[558],  nodes[353]);
    nmos (nodes[595], nodes[558],  nodes[354]);
    nmos (nodes[558], nodes[643],  nodes[444]);
    nmos (nodes[558], nodes[1613],  nodes[444]);
    nmos (nodes[1134], nodes[1431],  nodes[943]);
    nmos (nodes[256], nodes[558],  nodes[1478]);
    nmos (nodes[558], nodes[924],  nodes[1313]);
    nmos (nodes[710], nodes[558],  nodes[1105]);
    nmos (nodes[710], nodes[558],  nodes[1105]);
    nmos (nodes[558], nodes[710],  nodes[1105]);
    nmos (nodes[710], nodes[558],  nodes[1105]);
    nmos (nodes[558], nodes[710],  nodes[1105]);
    nmos (nodes[545], nodes[558],  nodes[1488]);
    nmos (nodes[1547], nodes[558],  nodes[1488]);
    nmos (nodes[815], nodes[558],  nodes[45]);
    nmos (nodes[570], nodes[558],  nodes[647]);
    nmos (nodes[1287], nodes[1491],  nodes[801]);
    nmos (nodes[558], nodes[467],  nodes[470]);
    nmos (nodes[737], nodes[146],  nodes[943]);
    nmos (nodes[1531], nodes[1188],  nodes[801]);
    nmos (nodes[558], nodes[513],  nodes[885]);
    nmos (nodes[37], nodes[558],  nodes[353]);
    nmos (nodes[37], nodes[558],  nodes[353]);
    nmos (nodes[313], nodes[350],  nodes[96]);
    nmos (nodes[558], nodes[649],  nodes[96]);
    nmos (nodes[798], nodes[558],  nodes[288]);
    nmos (nodes[794], nodes[657],  nodes[288]);
    nmos (nodes[657], nodes[826],  nodes[1429]);
    nmos (nodes[558], nodes[625],  nodes[43]);
    nmos (nodes[34], nodes[558],  nodes[1532]);
    nmos (nodes[652], nodes[558],  nodes[751]);
    nmos (nodes[475], nodes[558],  nodes[1677]);
    nmos (nodes[999], nodes[657],  nodes[1677]);
    nmos (nodes[958], nodes[865],  nodes[943]);
    nmos (nodes[85], nodes[1405],  nodes[1186]);
    nmos (nodes[1188], nodes[1648],  nodes[1186]);
    nmos (nodes[1287], nodes[1],  nodes[1186]);
    nmos (nodes[1067], nodes[558],  nodes[582]);
    nmos (nodes[657], nodes[821],  nodes[582]);
    nmos (nodes[448], nodes[1336],  nodes[1186]);
    nmos (nodes[166], nodes[589],  nodes[1186]);
    nmos (nodes[263], nodes[558],  nodes[1629]);
    nmos (nodes[1502], nodes[558],  nodes[707]);
    nmos (nodes[654], nodes[558],  nodes[71]);
    nmos (nodes[1001], nodes[777],  nodes[1186]);
    nmos (nodes[558], nodes[1719],  nodes[858]);
    nmos (nodes[558], nodes[1717],  nodes[60]);
    nmos (nodes[945], nodes[657],  nodes[520]);
    nmos (nodes[945], nodes[657],  nodes[520]);
    nmos (nodes[558], nodes[253],  nodes[1104]);
    nmos (nodes[558], nodes[362],  nodes[1552]);
    nmos (nodes[558], nodes[797],  nodes[892]);
    nmos (nodes[558], nodes[678],  nodes[644]);
    nmos (nodes[558], nodes[854],  nodes[975]);
    nmos (nodes[803], nodes[558],  nodes[1084]);
    nmos (nodes[558], nodes[1314],  nodes[1084]);
    nmos (nodes[1494], nodes[1454],  nodes[1205]);
    nmos (nodes[558], nodes[260],  nodes[1205]);
    nmos (nodes[982], nodes[1689],  nodes[943]);
    nmos (nodes[657], nodes[1001],  nodes[943]);
    nmos (nodes[88], nodes[522],  nodes[943]);
    nmos (nodes[914], nodes[484],  nodes[1386]);
    nmos (nodes[558], nodes[307],  nodes[31]);
    nmos (nodes[558], nodes[1580],  nodes[1287]);
    nmos (nodes[558], nodes[1580],  nodes[1287]);
    nmos (nodes[558], nodes[435],  nodes[86]);
    nmos (nodes[435], nodes[558],  nodes[86]);
    nmos (nodes[435], nodes[558],  nodes[86]);
    nmos (nodes[435], nodes[558],  nodes[86]);
    nmos (nodes[248], nodes[1624],  nodes[710]);
    nmos (nodes[558], nodes[616],  nodes[286]);
    nmos (nodes[558], nodes[482],  nodes[803]);
    nmos (nodes[736], nodes[558],  nodes[210]);
    nmos (nodes[736], nodes[558],  nodes[210]);
    nmos (nodes[736], nodes[558],  nodes[210]);
    nmos (nodes[736], nodes[558],  nodes[210]);
    nmos (nodes[558], nodes[959],  nodes[294]);
    nmos (nodes[1592], nodes[558],  nodes[128]);
    nmos (nodes[42], nodes[558],  nodes[353]);
    nmos (nodes[42], nodes[558],  nodes[353]);
    nmos (nodes[1613], nodes[558],  nodes[353]);
    nmos (nodes[1165], nodes[558],  nodes[910]);
    nmos (nodes[989], nodes[658],  nodes[943]);
    nmos (nodes[558], nodes[1304],  nodes[673]);
    nmos (nodes[558], nodes[39],  nodes[15]);
    nmos (nodes[880], nodes[1514],  nodes[710]);
    nmos (nodes[558], nodes[549],  nodes[708]);
    nmos (nodes[1531], nodes[305],  nodes[943]);
    nmos (nodes[629], nodes[202],  nodes[480]);
    nmos (nodes[1606], nodes[472],  nodes[710]);
    nmos (nodes[90], nodes[44],  nodes[943]);
    nmos (nodes[229], nodes[558],  nodes[683]);
    nmos (nodes[558], nodes[1380],  nodes[1154]);
    nmos (nodes[347], nodes[558],  nodes[904]);
    nmos (nodes[608], nodes[559],  nodes[943]);
    nmos (nodes[373], nodes[558],  nodes[353]);
    nmos (nodes[373], nodes[558],  nodes[353]);
    nmos (nodes[1720], nodes[558],  nodes[353]);
    nmos (nodes[657], nodes[54],  nodes[943]);
    nmos (nodes[68], nodes[722],  nodes[943]);
    nmos (nodes[302], nodes[558],  nodes[409]);
    nmos (nodes[957], nodes[841],  nodes[362]);
    nmos (nodes[681], nodes[250],  nodes[362]);
    nmos (nodes[740], nodes[350],  nodes[362]);
    nmos (nodes[1063], nodes[1071],  nodes[362]);
    nmos (nodes[477], nodes[296],  nodes[362]);
    nmos (nodes[336], nodes[277],  nodes[362]);
    nmos (nodes[1318], nodes[722],  nodes[362]);
    nmos (nodes[875], nodes[469],  nodes[943]);
    nmos (nodes[558], nodes[844],  nodes[1664]);
    nmos (nodes[1287], nodes[573],  nodes[325]);
    nmos (nodes[450], nodes[1656],  nodes[613]);
    nmos (nodes[1159], nodes[558],  nodes[613]);
    nmos (nodes[493], nodes[657],  nodes[943]);
    nmos (nodes[1452], nodes[1481],  nodes[943]);
    nmos (nodes[808], nodes[560],  nodes[943]);
    nmos (nodes[558], nodes[1517],  nodes[572]);
    nmos (nodes[1525], nodes[1348],  nodes[693]);
    nmos (nodes[558], nodes[169],  nodes[139]);
    nmos (nodes[1421], nodes[558],  nodes[334]);
    nmos (nodes[558], nodes[643],  nodes[353]);
    nmos (nodes[558], nodes[643],  nodes[353]);
    nmos (nodes[558], nodes[46],  nodes[248]);
    nmos (nodes[1185], nodes[558],  nodes[1137]);
    nmos (nodes[412], nodes[558],  nodes[560]);
    nmos (nodes[558], nodes[274],  nodes[860]);
    nmos (nodes[85], nodes[436],  nodes[943]);
    nmos (nodes[1284], nodes[896],  nodes[943]);
    nmos (nodes[180], nodes[558],  nodes[1716]);
    nmos (nodes[558], nodes[588],  nodes[1349]);
    nmos (nodes[1370], nodes[558],  nodes[1045]);
    nmos (nodes[132], nodes[1321],  nodes[943]);
    nmos (nodes[1307], nodes[1254],  nodes[943]);
    nmos (nodes[558], nodes[1347],  nodes[550]);
    nmos (nodes[816], nodes[1137],  nodes[790]);
    nmos (nodes[697], nodes[250],  nodes[943]);
    nmos (nodes[864], nodes[825],  nodes[639]);
    nmos (nodes[1588], nodes[558],  nodes[175]);
    nmos (nodes[1417], nodes[558],  nodes[747]);
    nmos (nodes[1309], nodes[558],  nodes[1460]);
    nmos (nodes[558], nodes[201],  nodes[1174]);
    nmos (nodes[798], nodes[558],  nodes[353]);
    nmos (nodes[798], nodes[558],  nodes[353]);
    nmos (nodes[288], nodes[558],  nodes[353]);
    nmos (nodes[525], nodes[558],  nodes[943]);
    nmos (nodes[628], nodes[558],  nodes[943]);
    nmos (nodes[558], nodes[1470],  nodes[1111]);
    nmos (nodes[1614], nodes[558],  nodes[1111]);
    nmos (nodes[558], nodes[313],  nodes[1680]);
    nmos (nodes[558], nodes[649],  nodes[1680]);
    nmos (nodes[558], nodes[984],  nodes[956]);
    nmos (nodes[242], nodes[558],  nodes[1521]);
    nmos (nodes[1150], nodes[1148],  nodes[325]);
    nmos (nodes[504], nodes[137],  nodes[440]);
    nmos (nodes[558], nodes[1649],  nodes[1382]);
    nmos (nodes[558], nodes[300],  nodes[1382]);
    nmos (nodes[558], nodes[1433],  nodes[90]);
    nmos (nodes[256], nodes[558],  nodes[120]);
    nmos (nodes[185], nodes[1063],  nodes[1645]);
    nmos (nodes[558], nodes[404],  nodes[1645]);
    nmos (nodes[1352], nodes[558],  nodes[1258]);
    nmos (nodes[1169], nodes[558],  nodes[987]);
    nmos (nodes[531], nodes[558],  nodes[95]);
    nmos (nodes[1051], nodes[31],  nodes[943]);
    nmos (nodes[1149], nodes[1368],  nodes[710]);
    nmos (nodes[558], nodes[612],  nodes[1453]);
    nmos (nodes[558], nodes[1720],  nodes[1453]);
    nmos (nodes[113], nodes[558],  nodes[126]);
    nmos (nodes[558], nodes[1391],  nodes[750]);
    nmos (nodes[1610], nodes[558],  nodes[640]);
    nmos (nodes[532], nodes[558],  nodes[1217]);
    nmos (nodes[558], nodes[476],  nodes[43]);
    nmos (nodes[1213], nodes[558],  nodes[453]);
    nmos (nodes[558], nodes[620],  nodes[1371]);
    nmos (nodes[558], nodes[51],  nodes[439]);
    nmos (nodes[334], nodes[558],  nodes[1553]);
    nmos (nodes[605], nodes[558],  nodes[1002]);
    nmos (nodes[605], nodes[558],  nodes[1002]);
    nmos (nodes[558], nodes[1541],  nodes[1477]);
    nmos (nodes[1107], nodes[558],  nodes[1428]);
    nmos (nodes[604], nodes[558],  nodes[1428]);
    nmos (nodes[89], nodes[558],  nodes[558]);
    nmos (nodes[272], nodes[558],  nodes[646]);
    nmos (nodes[1293], nodes[558],  nodes[1174]);
    nmos (nodes[1455], nodes[558],  nodes[131]);
    nmos (nodes[558], nodes[1331],  nodes[800]);
    nmos (nodes[741], nodes[558],  nodes[1247]);
    nmos (nodes[1014], nodes[121],  nodes[1564]);
    nmos (nodes[1387], nodes[1630],  nodes[1564]);
    nmos (nodes[266], nodes[1037],  nodes[943]);
    nmos (nodes[650], nodes[657],  nodes[42]);
    nmos (nodes[650], nodes[657],  nodes[42]);
    nmos (nodes[973], nodes[558],  nodes[1702]);
    nmos (nodes[1119], nodes[558],  nodes[1471]);
    nmos (nodes[621], nodes[1586],  nodes[943]);
    nmos (nodes[1046], nodes[577],  nodes[710]);
    nmos (nodes[956], nodes[558],  nodes[476]);
    nmos (nodes[657], nodes[984],  nodes[476]);
    nmos (nodes[558], nodes[1244],  nodes[1562]);
    nmos (nodes[558], nodes[1351],  nodes[1562]);
    nmos (nodes[558], nodes[961],  nodes[1503]);
    nmos (nodes[226], nodes[1093],  nodes[710]);
    nmos (nodes[558], nodes[1358],  nodes[245]);
    nmos (nodes[558], nodes[14],  nodes[671]);
    nmos (nodes[1662], nodes[558],  nodes[1124]);
    nmos (nodes[1401], nodes[558],  nodes[1269]);
    nmos (nodes[1249], nodes[558],  nodes[1269]);
    nmos (nodes[1451], nodes[668],  nodes[821]);
    nmos (nodes[558], nodes[1593],  nodes[226]);
    nmos (nodes[558], nodes[196],  nodes[543]);
    nmos (nodes[1468], nodes[657],  nodes[543]);
    nmos (nodes[236], nodes[558],  nodes[1708]);
    nmos (nodes[657], nodes[1237],  nodes[475]);
    nmos (nodes[558], nodes[827],  nodes[1350]);
    nmos (nodes[1472], nodes[827],  nodes[710]);
    nmos (nodes[1581], nodes[1275],  nodes[710]);
    nmos (nodes[1133], nodes[558],  nodes[1626]);
    nmos (nodes[702], nodes[558],  nodes[1626]);
    nmos (nodes[1353], nodes[1128],  nodes[821]);
    nmos (nodes[1037], nodes[558],  nodes[1086]);
    nmos (nodes[1105], nodes[558],  nodes[1399]);
    nmos (nodes[972], nodes[558],  nodes[319]);
    nmos (nodes[425], nodes[558],  nodes[936]);
    nmos (nodes[1005], nodes[657],  nodes[1325]);
    nmos (nodes[657], nodes[1005],  nodes[1325]);
    nmos (nodes[611], nodes[558],  nodes[43]);
    nmos (nodes[1106], nodes[558],  nodes[245]);
    nmos (nodes[1350], nodes[50],  nodes[710]);
    nmos (nodes[558], nodes[36],  nodes[600]);
    nmos (nodes[1048], nodes[558],  nodes[1721]);
    nmos (nodes[935], nodes[1636],  nodes[710]);
    nmos (nodes[558], nodes[503],  nodes[1394]);
    nmos (nodes[280], nodes[1630],  nodes[1468]);
    nmos (nodes[3], nodes[1437],  nodes[1468]);
    nmos (nodes[998], nodes[684],  nodes[1468]);
    nmos (nodes[1389], nodes[1242],  nodes[1468]);
    nmos (nodes[558], nodes[1004],  nodes[1408]);
    nmos (nodes[558], nodes[553],  nodes[1662]);
    nmos (nodes[1299], nodes[721],  nodes[1468]);
    nmos (nodes[558], nodes[1347],  nodes[862]);
    nmos (nodes[376], nodes[558],  nodes[107]);
    nmos (nodes[1151], nodes[182],  nodes[236]);
    nmos (nodes[141], nodes[558],  nodes[124]);
    nmos (nodes[1215], nodes[1528],  nodes[710]);
    nmos (nodes[109], nodes[1161],  nodes[710]);
    nmos (nodes[1198], nodes[626],  nodes[1401]);
    nmos (nodes[391], nodes[558],  nodes[529]);
    nmos (nodes[391], nodes[558],  nodes[529]);
    nmos (nodes[391], nodes[558],  nodes[529]);
    nmos (nodes[19], nodes[558],  nodes[770]);
    nmos (nodes[657], nodes[1150],  nodes[943]);
    nmos (nodes[265], nodes[182],  nodes[943]);
    nmos (nodes[1211], nodes[897],  nodes[943]);
    nmos (nodes[558], nodes[368],  nodes[446]);
    nmos (nodes[1354], nodes[558],  nodes[1165]);
    nmos (nodes[879], nodes[558],  nodes[1214]);
    nmos (nodes[558], nodes[1635],  nodes[966]);
    nmos (nodes[203], nodes[657],  nodes[966]);
    nmos (nodes[558], nodes[770],  nodes[559]);
    nmos (nodes[558], nodes[1271],  nodes[1596]);
    nmos (nodes[140], nodes[657],  nodes[1596]);
    nmos (nodes[1242], nodes[657],  nodes[943]);
    nmos (nodes[114], nodes[1402],  nodes[943]);
    nmos (nodes[1116], nodes[1014],  nodes[710]);
    nmos (nodes[1495], nodes[1546],  nodes[1600]);
    nmos (nodes[558], nodes[1044],  nodes[31]);
    nmos (nodes[979], nodes[558],  nodes[905]);
    nmos (nodes[558], nodes[156],  nodes[1533]);
    nmos (nodes[175], nodes[657],  nodes[373]);
    nmos (nodes[175], nodes[657],  nodes[373]);
    nmos (nodes[267], nodes[558],  nodes[1175]);
    nmos (nodes[657], nodes[1473],  nodes[943]);
    nmos (nodes[558], nodes[882],  nodes[597]);
    nmos (nodes[558], nodes[1056],  nodes[761]);
    nmos (nodes[619], nodes[695],  nodes[78]);
    nmos (nodes[1179], nodes[558],  nodes[78]);
    nmos (nodes[745], nodes[674],  nodes[943]);
    nmos (nodes[512], nodes[1130],  nodes[943]);
    nmos (nodes[1099], nodes[1102],  nodes[943]);
    nmos (nodes[558], nodes[269],  nodes[1241]);
    nmos (nodes[298], nodes[558],  nodes[353]);
    nmos (nodes[298], nodes[558],  nodes[353]);
    nmos (nodes[23], nodes[558],  nodes[353]);
    nmos (nodes[558], nodes[1279],  nodes[600]);
    nmos (nodes[969], nodes[558],  nodes[161]);
    nmos (nodes[801], nodes[657],  nodes[161]);
    nmos (nodes[558], nodes[715],  nodes[641]);
    nmos (nodes[558], nodes[1704],  nodes[641]);
    nmos (nodes[654], nodes[558],  nodes[1247]);
    nmos (nodes[604], nodes[558],  nodes[804]);
    nmos (nodes[166], nodes[615],  nodes[325]);
    nmos (nodes[1042], nodes[558],  nodes[1577]);
    nmos (nodes[414], nodes[558],  nodes[1043]);
    nmos (nodes[1001], nodes[843],  nodes[325]);
    nmos (nodes[558], nodes[1257],  nodes[1218]);
    nmos (nodes[558], nodes[1587],  nodes[894]);
    nmos (nodes[490], nodes[558],  nodes[1393]);
    nmos (nodes[557], nodes[1073],  nodes[344]);
    nmos (nodes[230], nodes[657],  nodes[826]);
    nmos (nodes[585], nodes[20],  nodes[344]);
    nmos (nodes[1316], nodes[558],  nodes[344]);
    nmos (nodes[934], nodes[73],  nodes[943]);
    nmos (nodes[558], nodes[1465],  nodes[248]);
    nmos (nodes[558], nodes[1349],  nodes[1501]);
    nmos (nodes[558], nodes[1349],  nodes[1501]);
    nmos (nodes[1349], nodes[558],  nodes[1501]);
    nmos (nodes[558], nodes[1349],  nodes[1501]);
    nmos (nodes[160], nodes[1049],  nodes[943]);
    nmos (nodes[558], nodes[647],  nodes[477]);
    nmos (nodes[264], nodes[558],  nodes[1149]);
    nmos (nodes[1218], nodes[558],  nodes[1565]);
    nmos (nodes[1218], nodes[558],  nodes[1565]);
    nmos (nodes[1276], nodes[248],  nodes[710]);
    nmos (nodes[501], nodes[1713],  nodes[943]);
    nmos (nodes[558], nodes[1512],  nodes[971]);
    nmos (nodes[558], nodes[258],  nodes[971]);
    nmos (nodes[558], nodes[84],  nodes[971]);
    nmos (nodes[558], nodes[788],  nodes[971]);
    nmos (nodes[558], nodes[1057],  nodes[971]);
    nmos (nodes[558], nodes[204],  nodes[971]);
    nmos (nodes[558], nodes[1582],  nodes[971]);
    nmos (nodes[558], nodes[1204],  nodes[971]);
    nmos (nodes[558], nodes[712],  nodes[971]);
    nmos (nodes[558], nodes[157],  nodes[971]);
    nmos (nodes[558], nodes[1086],  nodes[971]);
    nmos (nodes[558], nodes[487],  nodes[971]);
    nmos (nodes[558], nodes[1239],  nodes[971]);
    nmos (nodes[558], nodes[285],  nodes[971]);
    nmos (nodes[558], nodes[1524],  nodes[971]);
    nmos (nodes[558], nodes[273],  nodes[971]);
    nmos (nodes[558], nodes[750],  nodes[971]);
    nmos (nodes[558], nodes[932],  nodes[971]);
    nmos (nodes[558], nodes[309],  nodes[971]);
    nmos (nodes[558], nodes[219],  nodes[971]);
    nmos (nodes[1091], nodes[1360],  nodes[710]);
    nmos (nodes[1106], nodes[558],  nodes[84]);
    nmos (nodes[1262], nodes[558],  nodes[1679]);
    nmos (nodes[504], nodes[1438],  nodes[943]);
    nmos (nodes[1574], nodes[1228],  nodes[943]);
    nmos (nodes[1640], nodes[558],  nodes[843]);
    nmos (nodes[702], nodes[119],  nodes[943]);
    nmos (nodes[558], nodes[1006],  nodes[328]);
    nmos (nodes[119], nodes[237],  nodes[879]);
    nmos (nodes[310], nodes[724],  nodes[879]);
    nmos (nodes[1272], nodes[248],  nodes[710]);
    nmos (nodes[270], nodes[558],  nodes[503]);
    nmos (nodes[558], nodes[1684],  nodes[833]);
    nmos (nodes[256], nodes[558],  nodes[0]);
    nmos (nodes[1303], nodes[508],  nodes[335]);
    nmos (nodes[558], nodes[1460],  nodes[1669]);
    nmos (nodes[452], nodes[681],  nodes[704]);
    nmos (nodes[558], nodes[1691],  nodes[704]);
    nmos (nodes[737], nodes[54],  nodes[534]);
    nmos (nodes[1234], nodes[1009],  nodes[534]);
    nmos (nodes[450], nodes[978],  nodes[534]);
    nmos (nodes[162], nodes[1475],  nodes[534]);
    nmos (nodes[727], nodes[1405],  nodes[534]);
    nmos (nodes[858], nodes[263],  nodes[534]);
    nmos (nodes[1136], nodes[679],  nodes[534]);
    nmos (nodes[1653], nodes[1494],  nodes[534]);
    nmos (nodes[1028], nodes[558],  nodes[251]);
    nmos (nodes[558], nodes[353],  nodes[251]);
    nmos (nodes[558], nodes[353],  nodes[251]);
    nmos (nodes[353], nodes[558],  nodes[251]);
    nmos (nodes[353], nodes[558],  nodes[251]);
    nmos (nodes[558], nodes[19],  nodes[1708]);
    nmos (nodes[1108], nodes[54],  nodes[1060]);
    nmos (nodes[991], nodes[1150],  nodes[1060]);
    nmos (nodes[1287], nodes[1473],  nodes[1060]);
    nmos (nodes[1302], nodes[1188],  nodes[1060]);
    nmos (nodes[1405], nodes[892],  nodes[1060]);
    nmos (nodes[166], nodes[1503],  nodes[1060]);
    nmos (nodes[1336], nodes[833],  nodes[1060]);
    nmos (nodes[493], nodes[1001],  nodes[1060]);
    nmos (nodes[1124], nodes[1065],  nodes[943]);
    nmos (nodes[558], nodes[1144],  nodes[1571]);
    nmos (nodes[439], nodes[558],  nodes[1194]);
    nmos (nodes[1178], nodes[558],  nodes[848]);
    nmos (nodes[398], nodes[824],  nodes[943]);
    nmos (nodes[558], nodes[728],  nodes[1465]);
    nmos (nodes[1372], nodes[972],  nodes[388]);
    nmos (nodes[1250], nodes[558],  nodes[825]);
    nmos (nodes[742], nodes[558],  nodes[943]);
    nmos (nodes[454], nodes[558],  nodes[616]);
    nmos (nodes[774], nodes[558],  nodes[1419]);
    nmos (nodes[558], nodes[1258],  nodes[390]);
    nmos (nodes[558], nodes[1415],  nodes[1418]);
    nmos (nodes[1299], nodes[1147],  nodes[1564]);
    nmos (nodes[922], nodes[558],  nodes[620]);
    nmos (nodes[558], nodes[1115],  nodes[620]);
    nmos (nodes[1238], nodes[558],  nodes[1295]);
    nmos (nodes[1060], nodes[657],  nodes[1295]);
    nmos (nodes[663], nodes[1209],  nodes[943]);
    nmos (nodes[69], nodes[1181],  nodes[710]);
    nmos (nodes[171], nodes[28],  nodes[943]);
    nmos (nodes[558], nodes[437],  nodes[1247]);
    nmos (nodes[558], nodes[252],  nodes[1710]);
    nmos (nodes[558], nodes[1339],  nodes[799]);
    nmos (nodes[650], nodes[558],  nodes[643]);
    nmos (nodes[650], nodes[558],  nodes[643]);
    nmos (nodes[650], nodes[558],  nodes[643]);
    nmos (nodes[558], nodes[650],  nodes[643]);
    nmos (nodes[558], nodes[650],  nodes[643]);
    nmos (nodes[650], nodes[558],  nodes[643]);
    nmos (nodes[650], nodes[558],  nodes[643]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[1156], nodes[657],  nodes[102]);
    nmos (nodes[592], nodes[558],  nodes[1314]);
    nmos (nodes[1617], nodes[1327],  nodes[1314]);
    nmos (nodes[558], nodes[302],  nodes[1083]);
    nmos (nodes[558], nodes[1019],  nodes[1083]);
    nmos (nodes[648], nodes[558],  nodes[1200]);
    nmos (nodes[558], nodes[548],  nodes[1435]);
    nmos (nodes[558], nodes[1277],  nodes[1020]);
    nmos (nodes[558], nodes[1723],  nodes[1436]);
    nmos (nodes[1614], nodes[558],  nodes[1436]);
    nmos (nodes[903], nodes[1631],  nodes[1184]);
    nmos (nodes[657], nodes[1651],  nodes[943]);
    nmos (nodes[1172], nodes[1085],  nodes[372]);
    nmos (nodes[1290], nodes[912],  nodes[248]);
    nmos (nodes[773], nodes[558],  nodes[273]);
    nmos (nodes[17], nodes[558],  nodes[964]);
    nmos (nodes[1536], nodes[558],  nodes[964]);
    nmos (nodes[535], nodes[558],  nodes[663]);
    nmos (nodes[558], nodes[1286],  nodes[470]);
    nmos (nodes[558], nodes[135],  nodes[127]);
    nmos (nodes[901], nodes[558],  nodes[872]);
    nmos (nodes[1723], nodes[299],  nodes[1245]);
    nmos (nodes[657], nodes[1340],  nodes[1152]);
    nmos (nodes[657], nodes[1340],  nodes[1152]);
    nmos (nodes[1340], nodes[657],  nodes[1152]);
    nmos (nodes[1340], nodes[657],  nodes[1152]);
    nmos (nodes[657], nodes[1340],  nodes[1152]);
    nmos (nodes[558], nodes[1081],  nodes[1560]);
    nmos (nodes[558], nodes[1329],  nodes[1609]);
    nmos (nodes[558], nodes[1499],  nodes[1450]);
    nmos (nodes[1712], nodes[558],  nodes[926]);
    nmos (nodes[566], nodes[661],  nodes[1170]);
    nmos (nodes[1073], nodes[1326],  nodes[943]);
    nmos (nodes[7], nodes[558],  nodes[466]);
    nmos (nodes[471], nodes[657],  nodes[466]);
    nmos (nodes[558], nodes[384],  nodes[1258]);
    nmos (nodes[558], nodes[22],  nodes[193]);
    nmos (nodes[558], nodes[997],  nodes[289]);
    nmos (nodes[521], nodes[1358],  nodes[943]);
    nmos (nodes[1444], nodes[558],  nodes[318]);
    nmos (nodes[657], nodes[1443],  nodes[1545]);
    nmos (nodes[428], nodes[644],  nodes[710]);
    nmos (nodes[519], nodes[558],  nodes[1171]);
    nmos (nodes[558], nodes[1089],  nodes[1574]);
    nmos (nodes[1219], nodes[558],  nodes[776]);
    nmos (nodes[558], nodes[184],  nodes[305]);
    nmos (nodes[558], nodes[1079],  nodes[1411]);
    nmos (nodes[247], nodes[558],  nodes[849]);
    nmos (nodes[558], nodes[1211],  nodes[862]);
    nmos (nodes[1024], nodes[558],  nodes[94]);
    nmos (nodes[877], nodes[558],  nodes[933]);
    nmos (nodes[1406], nodes[1657],  nodes[523]);
    nmos (nodes[1659], nodes[875],  nodes[523]);
    nmos (nodes[743], nodes[558],  nodes[523]);
    nmos (nodes[513], nodes[558],  nodes[1646]);
    nmos (nodes[558], nodes[708],  nodes[1230]);
    nmos (nodes[549], nodes[657],  nodes[1230]);
    nmos (nodes[1398], nodes[304],  nodes[59]);
    nmos (nodes[957], nodes[143],  nodes[59]);
    nmos (nodes[1654], nodes[558],  nodes[947]);
    nmos (nodes[232], nodes[558],  nodes[377]);
    nmos (nodes[332], nodes[413],  nodes[1468]);
    nmos (nodes[558], nodes[1622],  nodes[758]);
    nmos (nodes[1190], nodes[558],  nodes[81]);
    nmos (nodes[1182], nodes[1300],  nodes[943]);
    nmos (nodes[1544], nodes[922],  nodes[270]);
    nmos (nodes[558], nodes[1115],  nodes[270]);
    nmos (nodes[110], nodes[558],  nodes[1691]);
    nmos (nodes[1023], nodes[558],  nodes[1691]);
    nmos (nodes[558], nodes[723],  nodes[868]);
    nmos (nodes[558], nodes[794],  nodes[746]);
    nmos (nodes[558], nodes[288],  nodes[746]);
    nmos (nodes[558], nodes[1681],  nodes[546]);
    nmos (nodes[558], nodes[1270],  nodes[43]);
    nmos (nodes[558], nodes[898],  nodes[1247]);
    nmos (nodes[1626], nodes[558],  nodes[119]);
    nmos (nodes[1197], nodes[1390],  nodes[500]);
    nmos (nodes[174], nodes[558],  nodes[500]);
    nmos (nodes[558], nodes[690],  nodes[188]);
    nmos (nodes[1040], nodes[782],  nodes[1303]);
    nmos (nodes[558], nodes[212],  nodes[1160]);
    nmos (nodes[819], nodes[558],  nodes[449]);
    nmos (nodes[558], nodes[457],  nodes[1302]);
    nmos (nodes[1015], nodes[558],  nodes[1033]);
    nmos (nodes[1299], nodes[1611],  nodes[414]);
    nmos (nodes[1188], nodes[305],  nodes[325]);
    nmos (nodes[55], nodes[11],  nodes[943]);
    nmos (nodes[1069], nodes[558],  nodes[1274]);
    nmos (nodes[1274], nodes[913],  nodes[710]);
    nmos (nodes[604], nodes[558],  nodes[1311]);
    nmos (nodes[298], nodes[558],  nodes[23]);
    nmos (nodes[1501], nodes[657],  nodes[23]);
    nmos (nodes[558], nodes[1093],  nodes[968]);
    nmos (nodes[1020], nodes[1705],  nodes[943]);
    nmos (nodes[781], nodes[558],  nodes[199]);
    nmos (nodes[1422], nodes[558],  nodes[199]);
    nmos (nodes[118], nodes[558],  nodes[334]);
    nmos (nodes[558], nodes[619],  nodes[700]);
    nmos (nodes[1090], nodes[558],  nodes[157]);
    nmos (nodes[1467], nodes[558],  nodes[1129]);
    nmos (nodes[736], nodes[657],  nodes[1633]);
    nmos (nodes[736], nodes[657],  nodes[1633]);
    nmos (nodes[736], nodes[657],  nodes[1633]);
    nmos (nodes[736], nodes[657],  nodes[1633]);
    nmos (nodes[736], nodes[657],  nodes[1633]);
    nmos (nodes[558], nodes[1556],  nodes[901]);
    nmos (nodes[558], nodes[867],  nodes[901]);
    nmos (nodes[558], nodes[1220],  nodes[647]);
    nmos (nodes[558], nodes[821],  nodes[1067]);
    nmos (nodes[1320], nodes[541],  nodes[943]);
    nmos (nodes[916], nodes[1409],  nodes[710]);
    nmos (nodes[862], nodes[558],  nodes[666]);
    nmos (nodes[558], nodes[283],  nodes[1323]);
    nmos (nodes[1206], nodes[558],  nodes[535]);
    nmos (nodes[558], nodes[1215],  nodes[1185]);
    nmos (nodes[558], nodes[1433],  nodes[201]);
    nmos (nodes[558], nodes[1200],  nodes[493]);
    nmos (nodes[744], nodes[558],  nodes[493]);
    nmos (nodes[967], nodes[558],  nodes[636]);
    nmos (nodes[657], nodes[268],  nodes[855]);
    nmos (nodes[657], nodes[268],  nodes[855]);
    nmos (nodes[657], nodes[268],  nodes[855]);
    nmos (nodes[657], nodes[268],  nodes[855]);
    nmos (nodes[657], nodes[268],  nodes[855]);
    nmos (nodes[1343], nodes[558],  nodes[248]);
    nmos (nodes[558], nodes[202],  nodes[646]);
    nmos (nodes[881], nodes[558],  nodes[943]);
    nmos (nodes[739], nodes[1080],  nodes[1056]);
    nmos (nodes[657], nodes[1539],  nodes[943]);
    nmos (nodes[558], nodes[631],  nodes[878]);
    nmos (nodes[1185], nodes[558],  nodes[916]);
    nmos (nodes[272], nodes[558],  nodes[967]);
    nmos (nodes[1333], nodes[80],  nodes[943]);
    nmos (nodes[558], nodes[571],  nodes[1671]);
    nmos (nodes[302], nodes[558],  nodes[1671]);
    nmos (nodes[558], nodes[1019],  nodes[1671]);
    nmos (nodes[1294], nodes[558],  nodes[1671]);
    nmos (nodes[558], nodes[1306],  nodes[1516]);
    nmos (nodes[1306], nodes[558],  nodes[1516]);
    nmos (nodes[558], nodes[1306],  nodes[1516]);
    nmos (nodes[1468], nodes[558],  nodes[196]);
    nmos (nodes[1058], nodes[558],  nodes[271]);
    nmos (nodes[24], nodes[1039],  nodes[710]);
    nmos (nodes[1649], nodes[558],  nodes[857]);
    nmos (nodes[1377], nodes[558],  nodes[857]);
    nmos (nodes[190], nodes[1101],  nodes[943]);
    nmos (nodes[558], nodes[412],  nodes[164]);
    nmos (nodes[20], nodes[993],  nodes[943]);
    nmos (nodes[558], nodes[726],  nodes[0]);
    nmos (nodes[558], nodes[1412],  nodes[1455]);
    nmos (nodes[1296], nodes[558],  nodes[1346]);
    nmos (nodes[657], nodes[359],  nodes[1346]);
    nmos (nodes[1455], nodes[558],  nodes[1324]);
    nmos (nodes[1001], nodes[765],  nodes[214]);
    nmos (nodes[104], nodes[558],  nodes[847]);
    nmos (nodes[1455], nodes[558],  nodes[1243]);
    nmos (nodes[148], nodes[558],  nodes[676]);
    nmos (nodes[558], nodes[148],  nodes[676]);
    nmos (nodes[148], nodes[558],  nodes[676]);
    nmos (nodes[558], nodes[148],  nodes[676]);
    nmos (nodes[148], nodes[558],  nodes[676]);
    nmos (nodes[148], nodes[558],  nodes[676]);
    nmos (nodes[148], nodes[558],  nodes[676]);
    nmos (nodes[1241], nodes[558],  nodes[748]);
    nmos (nodes[657], nodes[399],  nodes[1296]);
    nmos (nodes[267], nodes[558],  nodes[785]);
    nmos (nodes[657], nodes[353],  nodes[1028]);
    nmos (nodes[450], nodes[558],  nodes[1159]);
    nmos (nodes[558], nodes[1578],  nodes[1431]);
    nmos (nodes[558], nodes[1215],  nodes[238]);
    nmos (nodes[558], nodes[801],  nodes[969]);
    nmos (nodes[585], nodes[558],  nodes[232]);
    nmos (nodes[558], nodes[1704],  nodes[232]);
    nmos (nodes[1316], nodes[558],  nodes[232]);
    nmos (nodes[1069], nodes[1177],  nodes[943]);
    nmos (nodes[558], nodes[1315],  nodes[1429]);
    nmos (nodes[558], nodes[381],  nodes[1429]);
    nmos (nodes[1045], nodes[1442],  nodes[943]);
    nmos (nodes[1134], nodes[558],  nodes[1481]);
    nmos (nodes[357], nodes[728],  nodes[943]);
    nmos (nodes[160], nodes[558],  nodes[781]);
    nmos (nodes[912], nodes[558],  nodes[1481]);
    nmos (nodes[385], nodes[1652],  nodes[943]);
    nmos (nodes[558], nodes[1005],  nodes[558]);
    nmos (nodes[558], nodes[470],  nodes[646]);
    nmos (nodes[99], nodes[1194],  nodes[943]);
    nmos (nodes[558], nodes[556],  nodes[727]);
    nmos (nodes[558], nodes[368],  nodes[932]);
    nmos (nodes[1352], nodes[558],  nodes[932]);
    nmos (nodes[558], nodes[291],  nodes[1121]);
    nmos (nodes[733], nodes[558],  nodes[981]);
    nmos (nodes[66], nodes[107],  nodes[943]);
    nmos (nodes[657], nodes[475],  nodes[1143]);
    nmos (nodes[1677], nodes[558],  nodes[1143]);
    nmos (nodes[999], nodes[558],  nodes[1143]);
    nmos (nodes[394], nodes[957],  nodes[943]);
    nmos (nodes[558], nodes[1506],  nodes[1285]);
    nmos (nodes[1122], nodes[1510],  nodes[1285]);
    nmos (nodes[1175], nodes[558],  nodes[1447]);
    nmos (nodes[558], nodes[808],  nodes[1327]);
    nmos (nodes[558], nodes[1154],  nodes[959]);
    nmos (nodes[1493], nodes[558],  nodes[171]);
    nmos (nodes[1493], nodes[558],  nodes[171]);
    nmos (nodes[1493], nodes[558],  nodes[171]);
    nmos (nodes[1493], nodes[558],  nodes[171]);
    nmos (nodes[1686], nodes[1475],  nodes[345]);
    nmos (nodes[1097], nodes[558],  nodes[345]);
    nmos (nodes[767], nodes[558],  nodes[1138]);
    nmos (nodes[240], nodes[1387],  nodes[710]);
    nmos (nodes[1193], nodes[558],  nodes[815]);
    nmos (nodes[1065], nodes[558],  nodes[1292]);
    nmos (nodes[558], nodes[667],  nodes[829]);
    nmos (nodes[558], nodes[1434],  nodes[98]);
    nmos (nodes[558], nodes[830],  nodes[1505]);
    nmos (nodes[558], nodes[1030],  nodes[757]);
    nmos (nodes[671], nodes[1718],  nodes[710]);
    nmos (nodes[558], nodes[1130],  nodes[192]);
    nmos (nodes[1069], nodes[558],  nodes[1024]);
    nmos (nodes[1176], nodes[1231],  nodes[943]);
    nmos (nodes[558], nodes[1429],  nodes[1062]);
    nmos (nodes[358], nodes[558],  nodes[1171]);
    nmos (nodes[1090], nodes[558],  nodes[1222]);
    nmos (nodes[1717], nodes[558],  nodes[382]);
    nmos (nodes[54], nodes[1216],  nodes[1186]);
    nmos (nodes[482], nodes[1459],  nodes[336]);
    nmos (nodes[558], nodes[159],  nodes[558]);
    nmos (nodes[221], nodes[558],  nodes[1579]);
    nmos (nodes[892], nodes[1119],  nodes[1042]);
    nmos (nodes[558], nodes[374],  nodes[1591]);
    nmos (nodes[1302], nodes[439],  nodes[1042]);
    nmos (nodes[833], nodes[77],  nodes[1042]);
    nmos (nodes[558], nodes[279],  nodes[507]);
    nmos (nodes[1082], nodes[186],  nodes[507]);
    nmos (nodes[1266], nodes[961],  nodes[710]);
    nmos (nodes[1486], nodes[558],  nodes[200]);
    nmos (nodes[1367], nodes[293],  nodes[200]);
    nmos (nodes[57], nodes[558],  nodes[200]);
    nmos (nodes[558], nodes[1501],  nodes[353]);
    nmos (nodes[558], nodes[1501],  nodes[353]);
    nmos (nodes[1509], nodes[952],  nodes[943]);
    nmos (nodes[558], nodes[97],  nodes[222]);
    nmos (nodes[558], nodes[1245],  nodes[938]);
    nmos (nodes[1644], nodes[558],  nodes[99]);
    nmos (nodes[558], nodes[1666],  nodes[108]);
    nmos (nodes[558], nodes[1446],  nodes[850]);
    nmos (nodes[558], nodes[430],  nodes[850]);
    nmos (nodes[1216], nodes[1169],  nodes[943]);
    nmos (nodes[529], nodes[588],  nodes[943]);
    nmos (nodes[657], nodes[483],  nodes[943]);
    nmos (nodes[657], nodes[121],  nodes[943]);
    nmos (nodes[14], nodes[558],  nodes[67]);
    nmos (nodes[297], nodes[558],  nodes[1032]);
    nmos (nodes[763], nodes[558],  nodes[1534]);
    nmos (nodes[657], nodes[1068],  nodes[1534]);
    nmos (nodes[558], nodes[1045],  nodes[69]);
    nmos (nodes[1322], nodes[1009],  nodes[36]);
    nmos (nodes[735], nodes[558],  nodes[36]);
    nmos (nodes[539], nodes[657],  nodes[417]);
    nmos (nodes[657], nodes[539],  nodes[417]);
    nmos (nodes[657], nodes[539],  nodes[417]);
    nmos (nodes[539], nodes[657],  nodes[417]);
    nmos (nodes[539], nodes[657],  nodes[417]);
    nmos (nodes[539], nodes[657],  nodes[417]);
    nmos (nodes[657], nodes[539],  nodes[417]);
    nmos (nodes[558], nodes[1211],  nodes[967]);
    nmos (nodes[558], nodes[1211],  nodes[967]);
    nmos (nodes[558], nodes[1211],  nodes[1286]);
    nmos (nodes[1612], nodes[558],  nodes[690]);
    nmos (nodes[804], nodes[558],  nodes[690]);
    nmos (nodes[558], nodes[1311],  nodes[690]);
    nmos (nodes[558], nodes[492],  nodes[690]);
    nmos (nodes[558], nodes[1259],  nodes[690]);
    nmos (nodes[354], nodes[558],  nodes[690]);
    nmos (nodes[341], nodes[558],  nodes[690]);
    nmos (nodes[461], nodes[558],  nodes[690]);
    nmos (nodes[352], nodes[558],  nodes[690]);
    nmos (nodes[1589], nodes[558],  nodes[690]);
    nmos (nodes[558], nodes[1569],  nodes[690]);
    nmos (nodes[558], nodes[281],  nodes[690]);
    nmos (nodes[710], nodes[657],  nodes[1399]);
    nmos (nodes[558], nodes[321],  nodes[398]);
    nmos (nodes[558], nodes[692],  nodes[43]);
    nmos (nodes[558], nodes[620],  nodes[1293]);
    nmos (nodes[558], nodes[1122],  nodes[936]);
    nmos (nodes[558], nodes[1194],  nodes[348]);
    nmos (nodes[558], nodes[988],  nodes[350]);
    nmos (nodes[875], nodes[558],  nodes[743]);
    nmos (nodes[609], nodes[545],  nodes[743]);
    nmos (nodes[1547], nodes[558],  nodes[743]);
    nmos (nodes[1694], nodes[558],  nodes[890]);
    nmos (nodes[1001], nodes[1539],  nodes[140]);
    nmos (nodes[13], nodes[1336],  nodes[140]);
    nmos (nodes[54], nodes[64],  nodes[325]);
    nmos (nodes[54], nodes[407],  nodes[140]);
    nmos (nodes[558], nodes[38],  nodes[710]);
    nmos (nodes[1247], nodes[558],  nodes[710]);
    nmos (nodes[558], nodes[882],  nodes[1252]);
    nmos (nodes[1405], nodes[1160],  nodes[140]);
    nmos (nodes[1188], nodes[315],  nodes[140]);
    nmos (nodes[1287], nodes[1651],  nodes[140]);
    nmos (nodes[970], nodes[233],  nodes[761]);
    nmos (nodes[762], nodes[558],  nodes[761]);
    nmos (nodes[1372], nodes[558],  nodes[1201]);
    nmos (nodes[1293], nodes[558],  nodes[840]);
    nmos (nodes[558], nodes[1439],  nodes[115]);
    nmos (nodes[1072], nodes[558],  nodes[97]);
    nmos (nodes[769], nodes[558],  nodes[97]);
    nmos (nodes[1170], nodes[558],  nodes[755]);
    nmos (nodes[102], nodes[657],  nodes[834]);
    nmos (nodes[558], nodes[129],  nodes[75]);
    nmos (nodes[558], nodes[1571],  nodes[142]);
    nmos (nodes[165], nodes[427],  nodes[142]);
    nmos (nodes[957], nodes[1628],  nodes[574]);
    nmos (nodes[250], nodes[841],  nodes[574]);
    nmos (nodes[740], nodes[681],  nodes[574]);
    nmos (nodes[1071], nodes[350],  nodes[574]);
    nmos (nodes[296], nodes[1063],  nodes[574]);
    nmos (nodes[477], nodes[277],  nodes[574]);
    nmos (nodes[722], nodes[336],  nodes[574]);
    nmos (nodes[1318], nodes[304],  nodes[574]);
    nmos (nodes[569], nodes[1205],  nodes[233]);
    nmos (nodes[657], nodes[1282],  nodes[943]);
    nmos (nodes[887], nodes[657],  nodes[1191]);
    nmos (nodes[887], nodes[657],  nodes[1191]);
    nmos (nodes[887], nodes[657],  nodes[1191]);
    nmos (nodes[887], nodes[657],  nodes[1191]);
    nmos (nodes[709], nodes[558],  nodes[1499]);
    nmos (nodes[1201], nodes[657],  nodes[1499]);
    nmos (nodes[558], nodes[929],  nodes[1549]);
    nmos (nodes[558], nodes[414],  nodes[943]);
    nmos (nodes[558], nodes[898],  nodes[943]);
    nmos (nodes[132], nodes[558],  nodes[31]);
    nmos (nodes[558], nodes[1583],  nodes[918]);
    nmos (nodes[112], nodes[558],  nodes[336]);
    nmos (nodes[558], nodes[1110],  nodes[756]);
    nmos (nodes[1108], nodes[146],  nodes[1331]);
    nmos (nodes[991], nodes[929],  nodes[1331]);
    nmos (nodes[1473], nodes[1618],  nodes[1331]);
    nmos (nodes[1302], nodes[1654],  nodes[1331]);
    nmos (nodes[1344], nodes[892],  nodes[1331]);
    nmos (nodes[1503], nodes[831],  nodes[1331]);
    nmos (nodes[833], nodes[326],  nodes[1331]);
    nmos (nodes[493], nodes[1592],  nodes[1331]);
    nmos (nodes[558], nodes[540],  nodes[369]);
    nmos (nodes[1685], nodes[1542],  nodes[1345]);
    nmos (nodes[558], nodes[1568],  nodes[1345]);
    nmos (nodes[558], nodes[795],  nodes[1649]);
    nmos (nodes[1533], nodes[1180],  nodes[710]);
    nmos (nodes[983], nodes[558],  nodes[1403]);
    nmos (nodes[580], nodes[558],  nodes[1268]);
    nmos (nodes[1545], nodes[657],  nodes[287]);
    nmos (nodes[1034], nodes[558],  nodes[287]);
    nmos (nodes[994], nodes[558],  nodes[287]);
    nmos (nodes[347], nodes[558],  nodes[219]);
    nmos (nodes[52], nodes[1150],  nodes[140]);
    nmos (nodes[1332], nodes[558],  nodes[984]);
    nmos (nodes[582], nodes[558],  nodes[610]);
    nmos (nodes[1001], nodes[1251],  nodes[801]);
    nmos (nodes[558], nodes[937],  nodes[1139]);
    nmos (nodes[526], nodes[1500],  nodes[943]);
    nmos (nodes[1405], nodes[658],  nodes[801]);
    nmos (nodes[558], nodes[603],  nodes[47]);
    nmos (nodes[1336], nodes[518],  nodes[801]);
    nmos (nodes[166], nodes[733],  nodes[801]);
    nmos (nodes[558], nodes[499],  nodes[49]);
    nmos (nodes[824], nodes[558],  nodes[579]);
    nmos (nodes[445], nodes[558],  nodes[862]);
    nmos (nodes[1185], nodes[558],  nodes[729]);
    nmos (nodes[1519], nodes[738],  nodes[710]);
    nmos (nodes[734], nodes[558],  nodes[1540]);
    nmos (nodes[657], nodes[1503],  nodes[943]);
    nmos (nodes[629], nodes[558],  nodes[50]);
    nmos (nodes[151], nodes[440],  nodes[943]);
    nmos (nodes[558], nodes[1716],  nodes[660]);
    nmos (nodes[558], nodes[1708],  nodes[660]);
    nmos (nodes[256], nodes[558],  nodes[594]);
    nmos (nodes[208], nodes[558],  nodes[39]);
    nmos (nodes[1349], nodes[558],  nodes[558]);
    nmos (nodes[26], nodes[927],  nodes[943]);
    nmos (nodes[558], nodes[1335],  nodes[628]);
    nmos (nodes[1698], nodes[657],  nodes[628]);
    nmos (nodes[460], nodes[616],  nodes[943]);
    nmos (nodes[1233], nodes[558],  nodes[895]);
    nmos (nodes[76], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[1658],  nodes[895]);
    nmos (nodes[786], nodes[558],  nodes[895]);
    nmos (nodes[1664], nodes[558],  nodes[895]);
    nmos (nodes[1612], nodes[558],  nodes[895]);
    nmos (nodes[784], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[244],  nodes[895]);
    nmos (nodes[558], nodes[1623],  nodes[895]);
    nmos (nodes[764], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[1311],  nodes[895]);
    nmos (nodes[558], nodes[324],  nodes[895]);
    nmos (nodes[558], nodes[857],  nodes[895]);
    nmos (nodes[1337], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[1355],  nodes[895]);
    nmos (nodes[558], nodes[787],  nodes[895]);
    nmos (nodes[575], nodes[558],  nodes[895]);
    nmos (nodes[1381], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[822],  nodes[895]);
    nmos (nodes[558], nodes[131],  nodes[895]);
    nmos (nodes[1086], nodes[558],  nodes[895]);
    nmos (nodes[1074], nodes[558],  nodes[895]);
    nmos (nodes[1246], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[0],  nodes[895]);
    nmos (nodes[594], nodes[558],  nodes[895]);
    nmos (nodes[1052], nodes[558],  nodes[895]);
    nmos (nodes[1589], nodes[558],  nodes[895]);
    nmos (nodes[446], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[309],  nodes[895]);
    nmos (nodes[558], nodes[53],  nodes[895]);
    nmos (nodes[558], nodes[1292],  nodes[895]);
    nmos (nodes[1155], nodes[558],  nodes[895]);
    nmos (nodes[1569], nodes[558],  nodes[895]);
    nmos (nodes[301], nodes[558],  nodes[895]);
    nmos (nodes[950], nodes[558],  nodes[895]);
    nmos (nodes[1710], nodes[558],  nodes[895]);
    nmos (nodes[558], nodes[1419],  nodes[895]);
    nmos (nodes[716], nodes[558],  nodes[681]);
    nmos (nodes[1503], nodes[72],  nodes[283]);
    nmos (nodes[558], nodes[693],  nodes[143]);
    nmos (nodes[558], nodes[1285],  nodes[143]);
    nmos (nodes[604], nodes[558],  nodes[1031]);
    nmos (nodes[1505], nodes[1455],  nodes[943]);
    nmos (nodes[558], nodes[1240],  nodes[1566]);
    nmos (nodes[863], nodes[657],  nodes[1566]);
    nmos (nodes[864], nodes[1507],  nodes[710]);
    nmos (nodes[558], nodes[996],  nodes[1133]);
    nmos (nodes[919], nodes[856],  nodes[1704]);
    nmos (nodes[558], nodes[835],  nodes[1704]);
    nmos (nodes[558], nodes[838],  nodes[581]);
    nmos (nodes[1563], nodes[11],  nodes[397]);
    nmos (nodes[558], nodes[134],  nodes[1557]);
    nmos (nodes[208], nodes[892],  nodes[283]);
    nmos (nodes[558], nodes[1130],  nodes[862]);
    nmos (nodes[315], nodes[657],  nodes[943]);
    nmos (nodes[558], nodes[133],  nodes[943]);
    nmos (nodes[558], nodes[161],  nodes[943]);
    nmos (nodes[332], nodes[558],  nodes[418]);
    nmos (nodes[276], nodes[740],  nodes[943]);
    nmos (nodes[1000], nodes[558],  nodes[1466]);
    nmos (nodes[558], nodes[753],  nodes[1257]);
    nmos (nodes[558], nodes[711],  nodes[1257]);
    nmos (nodes[569], nodes[558],  nodes[1257]);
    nmos (nodes[558], nodes[440],  nodes[24]);
    nmos (nodes[558], nodes[1025],  nodes[64]);
    nmos (nodes[1107], nodes[558],  nodes[58]);
    nmos (nodes[360], nodes[795],  nodes[943]);
    nmos (nodes[1554], nodes[679],  nodes[739]);
    nmos (nodes[479], nodes[558],  nodes[739]);
    nmos (nodes[1631], nodes[868],  nodes[943]);
    nmos (nodes[272], nodes[558],  nodes[0]);
    nmos (nodes[1349], nodes[657],  nodes[298]);
    nmos (nodes[1349], nodes[657],  nodes[298]);
    nmos (nodes[1349], nodes[657],  nodes[298]);
    nmos (nodes[1349], nodes[657],  nodes[298]);
    nmos (nodes[195], nodes[558],  nodes[659]);
    nmos (nodes[558], nodes[195],  nodes[659]);
    nmos (nodes[558], nodes[195],  nodes[659]);
    nmos (nodes[558], nodes[195],  nodes[659]);
    nmos (nodes[195], nodes[558],  nodes[659]);
    nmos (nodes[558], nodes[195],  nodes[659]);
    nmos (nodes[146], nodes[54],  nodes[1698]);
    nmos (nodes[929], nodes[1150],  nodes[1698]);
    nmos (nodes[1287], nodes[1618],  nodes[1698]);
    nmos (nodes[1654], nodes[1188],  nodes[1698]);
    nmos (nodes[1344], nodes[1405],  nodes[1698]);
    nmos (nodes[831], nodes[166],  nodes[1698]);
    nmos (nodes[1336], nodes[326],  nodes[1698]);
    nmos (nodes[1001], nodes[1592],  nodes[1698]);
    nmos (nodes[694], nodes[1282],  nodes[1468]);
    nmos (nodes[642], nodes[707],  nodes[943]);
    nmos (nodes[558], nodes[1722],  nodes[780]);
    nmos (nodes[1704], nodes[558],  nodes[379]);
    nmos (nodes[558], nodes[1512],  nodes[1125]);
    nmos (nodes[382], nodes[558],  nodes[1125]);
    nmos (nodes[558], nodes[1173],  nodes[1125]);
    nmos (nodes[558], nodes[1543],  nodes[1125]);
    nmos (nodes[558], nodes[76],  nodes[1125]);
    nmos (nodes[558], nodes[245],  nodes[1125]);
    nmos (nodes[558], nodes[786],  nodes[1125]);
    nmos (nodes[558], nodes[1664],  nodes[1125]);
    nmos (nodes[558], nodes[682],  nodes[1125]);
    nmos (nodes[558], nodes[1482],  nodes[1125]);
    nmos (nodes[558], nodes[552],  nodes[1125]);
    nmos (nodes[558], nodes[1487],  nodes[1125]);
    nmos (nodes[558], nodes[764],  nodes[1125]);
    nmos (nodes[558], nodes[1057],  nodes[1125]);
    nmos (nodes[558], nodes[58],  nodes[1125]);
    nmos (nodes[558], nodes[1520],  nodes[1125]);
    nmos (nodes[558], nodes[1381],  nodes[1125]);
    nmos (nodes[558], nodes[257],  nodes[1125]);
    nmos (nodes[558], nodes[1324],  nodes[1125]);
    nmos (nodes[558], nodes[179],  nodes[1125]);
    nmos (nodes[131], nodes[558],  nodes[1125]);
    nmos (nodes[558], nodes[4],  nodes[1125]);
    nmos (nodes[558], nodes[1396],  nodes[1125]);
    nmos (nodes[558], nodes[167],  nodes[1125]);
    nmos (nodes[558], nodes[354],  nodes[1125]);
    nmos (nodes[558], nodes[1086],  nodes[1125]);
    nmos (nodes[558], nodes[1074],  nodes[1125]);
    nmos (nodes[273], nodes[558],  nodes[1125]);
    nmos (nodes[558], nodes[594],  nodes[1125]);
    nmos (nodes[558], nodes[677],  nodes[1125]);
    nmos (nodes[558], nodes[447],  nodes[1125]);
    nmos (nodes[558], nodes[1052],  nodes[1125]);
    nmos (nodes[791], nodes[558],  nodes[1125]);
    nmos (nodes[558], nodes[750],  nodes[1125]);
    nmos (nodes[558], nodes[932],  nodes[1125]);
    nmos (nodes[558], nodes[1589],  nodes[1125]);
    nmos (nodes[558], nodes[309],  nodes[1125]);
    nmos (nodes[558], nodes[1430],  nodes[1125]);
    nmos (nodes[558], nodes[1292],  nodes[1125]);
    nmos (nodes[558], nodes[1114],  nodes[1125]);
    nmos (nodes[558], nodes[1226],  nodes[1125]);
    nmos (nodes[558], nodes[1006],  nodes[1125]);
    nmos (nodes[558], nodes[1164],  nodes[1125]);
    nmos (nodes[558], nodes[950],  nodes[1125]);
    nmos (nodes[558], nodes[281],  nodes[1125]);
    nmos (nodes[558], nodes[1665],  nodes[1125]);
    nmos (nodes[558], nodes[607],  nodes[1125]);
    nmos (nodes[558], nodes[1419],  nodes[1125]);
    nmos (nodes[558], nodes[1050],  nodes[1125]);
    nmos (nodes[558], nodes[59],  nodes[1255]);
    nmos (nodes[558], nodes[1546],  nodes[781]);
    nmos (nodes[1457], nodes[558],  nodes[781]);
    nmos (nodes[1369], nodes[558],  nodes[897]);
    nmos (nodes[558], nodes[1508],  nodes[46]);
    nmos (nodes[1559], nodes[558],  nodes[530]);
    nmos (nodes[1632], nodes[558],  nodes[530]);
    nmos (nodes[510], nodes[558],  nodes[434]);
    nmos (nodes[558], nodes[414],  nodes[1247]);
    nmos (nodes[558], nodes[152],  nodes[630]);
    nmos (nodes[1572], nodes[558],  nodes[701]);
    nmos (nodes[193], nodes[558],  nodes[701]);
    nmos (nodes[558], nodes[1352],  nodes[335]);
    nmos (nodes[1156], nodes[558],  nodes[1696]);
    nmos (nodes[558], nodes[1156],  nodes[1696]);
    nmos (nodes[558], nodes[1156],  nodes[1696]);
    nmos (nodes[1156], nodes[558],  nodes[1696]);
    nmos (nodes[558], nodes[1156],  nodes[1696]);
    nmos (nodes[558], nodes[407],  nodes[229]);
    nmos (nodes[558], nodes[506],  nodes[192]);
    nmos (nodes[558], nodes[925],  nodes[517]);
    nmos (nodes[558], nodes[139],  nodes[934]);
    nmos (nodes[1711], nodes[1064],  nodes[943]);
    nmos (nodes[1443], nodes[657],  nodes[1545]);
    nmos (nodes[1181], nodes[648],  nodes[754]);
    nmos (nodes[558], nodes[1595],  nodes[754]);
    nmos (nodes[52], nodes[292],  nodes[48]);
    nmos (nodes[1178], nodes[590],  nodes[710]);
    nmos (nodes[775], nodes[558],  nodes[1128]);
    nmos (nodes[407], nodes[1670],  nodes[48]);
    nmos (nodes[558], nodes[617],  nodes[713]);
    nmos (nodes[558], nodes[676],  nodes[713]);
    nmos (nodes[1192], nodes[751],  nodes[943]);
    nmos (nodes[1639], nodes[657],  nodes[489]);
    nmos (nodes[1153], nodes[558],  nodes[489]);
    nmos (nodes[558], nodes[659],  nodes[489]);
    nmos (nodes[100], nodes[558],  nodes[1018]);
    nmos (nodes[558], nodes[1469],  nodes[1220]);
    nmos (nodes[778], nodes[558],  nodes[231]);
    nmos (nodes[368], nodes[558],  nodes[1430]);
    nmos (nodes[558], nodes[911],  nodes[877]);
    nmos (nodes[558], nodes[911],  nodes[877]);
    nmos (nodes[847], nodes[558],  nodes[300]);
    nmos (nodes[602], nodes[558],  nodes[133]);
    nmos (nodes[1263], nodes[657],  nodes[133]);
    nmos (nodes[558], nodes[1201],  nodes[709]);
    nmos (nodes[558], nodes[987],  nodes[1216]);
    nmos (nodes[1293], nodes[558],  nodes[318]);
    nmos (nodes[1075], nodes[558],  nodes[1393]);
    nmos (nodes[1007], nodes[558],  nodes[1704]);
    nmos (nodes[558], nodes[176],  nodes[236]);
    nmos (nodes[652], nodes[1551],  nodes[741]);
    nmos (nodes[1206], nodes[205],  nodes[741]);
    nmos (nodes[27], nodes[948],  nodes[741]);
    nmos (nodes[1301], nodes[49],  nodes[741]);
    nmos (nodes[1496], nodes[502],  nodes[741]);
    nmos (nodes[141], nodes[584],  nodes[741]);
    nmos (nodes[1722], nodes[1670],  nodes[741]);
    nmos (nodes[209], nodes[292],  nodes[741]);
    nmos (nodes[1411], nodes[515],  nodes[943]);
    nmos (nodes[558], nodes[616],  nodes[665]);
    nmos (nodes[315], nodes[558],  nodes[203]);
    nmos (nodes[1651], nodes[558],  nodes[203]);
    nmos (nodes[483], nodes[558],  nodes[203]);
    nmos (nodes[1160], nodes[558],  nodes[203]);
    nmos (nodes[558], nodes[550],  nodes[1228]);
    nmos (nodes[1539], nodes[558],  nodes[203]);
    nmos (nodes[13], nodes[558],  nodes[203]);
    nmos (nodes[558], nodes[1230],  nodes[360]);
    nmos (nodes[558], nodes[1118],  nodes[204]);
    nmos (nodes[1058], nodes[632],  nodes[1289]);
    nmos (nodes[198], nodes[558],  nodes[197]);
    nmos (nodes[198], nodes[558],  nodes[197]);
    nmos (nodes[1092], nodes[558],  nodes[888]);
    nmos (nodes[74], nodes[1675],  nodes[879]);
    nmos (nodes[1378], nodes[1609],  nodes[879]);
    nmos (nodes[1082], nodes[1692],  nodes[270]);
    nmos (nodes[558], nodes[1668],  nodes[407]);
    nmos (nodes[824], nodes[558],  nodes[487]);
    nmos (nodes[583], nodes[1432],  nodes[1068]);
    nmos (nodes[1621], nodes[96],  nodes[1068]);
    nmos (nodes[558], nodes[1619],  nodes[182]);
    nmos (nodes[1486], nodes[126],  nodes[943]);
    nmos (nodes[558], nodes[152],  nodes[788]);
    nmos (nodes[1492], nodes[558],  nodes[974]);
    nmos (nodes[558], nodes[378],  nodes[1357]);
    nmos (nodes[558], nodes[732],  nodes[1161]);
    nmos (nodes[1621], nodes[558],  nodes[1302]);
    nmos (nodes[182], nodes[558],  nodes[646]);
    nmos (nodes[347], nodes[558],  nodes[607]);
    nmos (nodes[1298], nodes[1267],  nodes[710]);
    nmos (nodes[42], nodes[558],  nodes[1613]);
    nmos (nodes[643], nodes[657],  nodes[1613]);
    nmos (nodes[1682], nodes[558],  nodes[901]);
    nmos (nodes[1362], nodes[558],  nodes[901]);
    nmos (nodes[378], nodes[940],  nodes[943]);
    nmos (nodes[187], nodes[558],  nodes[248]);
    nmos (nodes[1718], nodes[558],  nodes[248]);
    nmos (nodes[837], nodes[558],  nodes[1623]);
    nmos (nodes[657], nodes[1163],  nodes[747]);
    nmos (nodes[1715], nodes[558],  nodes[358]);
    nmos (nodes[208], nodes[1437],  nodes[438]);
    nmos (nodes[1630], nodes[72],  nodes[438]);
    nmos (nodes[1458], nodes[121],  nodes[438]);
    nmos (nodes[1299], nodes[1647],  nodes[438]);
    nmos (nodes[488], nodes[413],  nodes[438]);
    nmos (nodes[1282], nodes[976],  nodes[438]);
    nmos (nodes[481], nodes[1242],  nodes[438]);
    nmos (nodes[684], nodes[723],  nodes[438]);
    nmos (nodes[558], nodes[975],  nodes[854]);
    nmos (nodes[1500], nodes[558],  nodes[1345]);
    nmos (nodes[289], nodes[635],  nodes[943]);
    nmos (nodes[133], nodes[558],  nodes[1404]);
    nmos (nodes[1242], nodes[558],  nodes[1193]);
    nmos (nodes[1416], nodes[558],  nodes[833]);
    nmos (nodes[558], nodes[930],  nodes[1276]);
    nmos (nodes[558], nodes[930],  nodes[1276]);
    nmos (nodes[83], nodes[558],  nodes[1400]);
    nmos (nodes[558], nodes[611],  nodes[1509]);
    nmos (nodes[1507], nodes[558],  nodes[684]);
    nmos (nodes[657], nodes[43],  nodes[839]);
    nmos (nodes[536], nodes[484],  nodes[943]);
    nmos (nodes[558], nodes[6],  nodes[43]);
    nmos (nodes[1206], nodes[1539],  nodes[1235]);
    nmos (nodes[652], nodes[13],  nodes[1235]);
    nmos (nodes[1301], nodes[483],  nodes[1235]);
    nmos (nodes[27], nodes[1160],  nodes[1235]);
    nmos (nodes[141], nodes[315],  nodes[1235]);
    nmos (nodes[1496], nodes[1651],  nodes[1235]);
    nmos (nodes[209], nodes[52],  nodes[1235]);
    nmos (nodes[1722], nodes[407],  nodes[1235]);
    nmos (nodes[779], nodes[605],  nodes[1440]);
    nmos (nodes[700], nodes[558],  nodes[1201]);
    nmos (nodes[381], nodes[1062],  nodes[943]);
    nmos (nodes[558], nodes[1129],  nodes[710]);
    nmos (nodes[1352], nodes[558],  nodes[1642]);
    nmos (nodes[657], nodes[211],  nodes[1041]);
    nmos (nodes[211], nodes[657],  nodes[1041]);
    nmos (nodes[211], nodes[657],  nodes[1041]);
    nmos (nodes[211], nodes[657],  nodes[1041]);
    nmos (nodes[657], nodes[211],  nodes[1041]);
    nmos (nodes[558], nodes[1254],  nodes[178]);
    nmos (nodes[558], nodes[1195],  nodes[178]);
    nmos (nodes[1191], nodes[657],  nodes[178]);
    nmos (nodes[558], nodes[300],  nodes[389]);
    nmos (nodes[491], nodes[558],  nodes[1541]);
    nmos (nodes[657], nodes[437],  nodes[1541]);
    nmos (nodes[431], nodes[558],  nodes[943]);
    nmos (nodes[195], nodes[657],  nodes[1639]);
    nmos (nodes[657], nodes[1237],  nodes[475]);
    nmos (nodes[1072], nodes[558],  nodes[353]);
    nmos (nodes[1072], nodes[558],  nodes[353]);
    nmos (nodes[558], nodes[1189],  nodes[1008]);
    nmos (nodes[1511], nodes[558],  nodes[1008]);
    nmos (nodes[814], nodes[344],  nodes[410]);
    nmos (nodes[558], nodes[557],  nodes[410]);
    nmos (nodes[375], nodes[558],  nodes[308]);
    nmos (nodes[65], nodes[558],  nodes[308]);
    nmos (nodes[678], nodes[706],  nodes[943]);
    nmos (nodes[533], nodes[558],  nodes[561]);
    nmos (nodes[474], nodes[558],  nodes[410]);
    nmos (nodes[1608], nodes[558],  nodes[1423]);
    nmos (nodes[657], nodes[869],  nodes[1423]);
    nmos (nodes[836], nodes[168],  nodes[710]);
    nmos (nodes[558], nodes[1392],  nodes[1297]);
    nmos (nodes[1024], nodes[1699],  nodes[943]);
    nmos (nodes[1232], nodes[558],  nodes[364]);
    nmos (nodes[18], nodes[468],  nodes[710]);
    nmos (nodes[296], nodes[404],  nodes[59]);
    nmos (nodes[558], nodes[1649],  nodes[389]);
    nmos (nodes[1464], nodes[558],  nodes[1487]);
    nmos (nodes[277], nodes[1632],  nodes[59]);
    nmos (nodes[378], nodes[558],  nodes[18]);
    nmos (nodes[379], nodes[1480],  nodes[1570]);
    nmos (nodes[657], nodes[833],  nodes[943]);
    nmos (nodes[905], nodes[1681],  nodes[440]);
    nmos (nodes[576], nodes[213],  nodes[943]);
    nmos (nodes[537], nodes[862],  nodes[943]);
    nmos (nodes[158], nodes[789],  nodes[710]);
    nmos (nodes[558], nodes[1685],  nodes[1166]);
    nmos (nodes[558], nodes[1568],  nodes[1166]);
    nmos (nodes[855], nodes[558],  nodes[1660]);
    nmos (nodes[657], nodes[1100],  nodes[1660]);
    nmos (nodes[1712], nodes[558],  nodes[1134]);
    nmos (nodes[558], nodes[1006],  nodes[1050]);
    nmos (nodes[1594], nodes[656],  nodes[779]);
    nmos (nodes[1032], nodes[558],  nodes[297]);
    nmos (nodes[1344], nodes[558],  nodes[556]);
    nmos (nodes[1196], nodes[558],  nodes[1689]);
    nmos (nodes[826], nodes[558],  nodes[1315]);
    nmos (nodes[558], nodes[1202],  nodes[1265]);
    nmos (nodes[558], nodes[1334],  nodes[1265]);
    nmos (nodes[615], nodes[733],  nodes[943]);
    nmos (nodes[195], nodes[657],  nodes[1639]);
    nmos (nodes[558], nodes[63],  nodes[158]);
    nmos (nodes[1703], nodes[558],  nodes[1373]);
    nmos (nodes[395], nodes[558],  nodes[1373]);
    nmos (nodes[1639], nodes[558],  nodes[1153]);
    nmos (nodes[657], nodes[659],  nodes[1153]);
    nmos (nodes[558], nodes[761],  nodes[314]);
    nmos (nodes[1550], nodes[558],  nodes[781]);
    nmos (nodes[1269], nodes[967],  nodes[943]);
    nmos (nodes[1390], nodes[558],  nodes[1459]);
    nmos (nodes[174], nodes[558],  nodes[1459]);
    nmos (nodes[11], nodes[558],  nodes[1396]);
    nmos (nodes[327], nodes[199],  nodes[943]);
    nmos (nodes[338], nodes[252],  nodes[943]);
    nmos (nodes[1579], nodes[187],  nodes[710]);
    nmos (nodes[566], nodes[627],  nodes[710]);
    nmos (nodes[558], nodes[1186],  nodes[1247]);
    nmos (nodes[581], nodes[306],  nodes[943]);
    nmos (nodes[558], nodes[1564],  nodes[1157]);
    nmos (nodes[1374], nodes[558],  nodes[562]);
    nmos (nodes[558], nodes[1453],  nodes[1266]);
    nmos (nodes[657], nodes[195],  nodes[1639]);
    nmos (nodes[558], nodes[744],  nodes[1473]);
    nmos (nodes[314], nodes[558],  nodes[893]);
    nmos (nodes[1573], nodes[558],  nodes[1473]);
    nmos (nodes[558], nodes[662],  nodes[625]);
    nmos (nodes[1186], nodes[657],  nodes[625]);
    nmos (nodes[1172], nodes[558],  nodes[646]);
    nmos (nodes[464], nodes[558],  nodes[1284]);
    nmos (nodes[464], nodes[558],  nodes[1284]);
    nmos (nodes[464], nodes[558],  nodes[1284]);
    nmos (nodes[505], nodes[558],  nodes[1122]);
    nmos (nodes[433], nodes[558],  nodes[1122]);
    nmos (nodes[1213], nodes[558],  nodes[609]);
    nmos (nodes[657], nodes[1325],  nodes[97]);
    nmos (nodes[385], nodes[558],  nodes[604]);
    nmos (nodes[558], nodes[522],  nodes[1145]);
    nmos (nodes[5], nodes[558],  nodes[737]);
    nmos (nodes[1717], nodes[558],  nodes[1512]);
    nmos (nodes[17], nodes[554],  nodes[943]);
    nmos (nodes[1615], nodes[558],  nodes[940]);
    nmos (nodes[558], nodes[399],  nodes[359]);
    nmos (nodes[558], nodes[399],  nodes[359]);
    nmos (nodes[399], nodes[558],  nodes[359]);
    nmos (nodes[558], nodes[399],  nodes[359]);
    nmos (nodes[399], nodes[558],  nodes[359]);
    nmos (nodes[558], nodes[399],  nodes[359]);
    nmos (nodes[558], nodes[399],  nodes[359]);
    nmos (nodes[558], nodes[191],  nodes[790]);
    nmos (nodes[558], nodes[1107],  nodes[1204]);
    nmos (nodes[1638], nodes[558],  nodes[1591]);
    nmos (nodes[836], nodes[768],  nodes[821]);
    nmos (nodes[465], nodes[558],  nodes[206]);
    nmos (nodes[368], nodes[558],  nodes[528]);
    nmos (nodes[558], nodes[316],  nodes[1167]);
    nmos (nodes[143], nodes[558],  nodes[1167]);
    nmos (nodes[558], nodes[696],  nodes[217]);
    nmos (nodes[558], nodes[210],  nodes[234]);
    nmos (nodes[558], nodes[172],  nodes[234]);
    nmos (nodes[657], nodes[1633],  nodes[234]);
    nmos (nodes[558], nodes[1618],  nodes[419]);
    nmos (nodes[558], nodes[43],  nodes[710]);
    nmos (nodes[1247], nodes[558],  nodes[710]);
    nmos (nodes[558], nodes[1247],  nodes[710]);
    nmos (nodes[947], nodes[558],  nodes[162]);
    nmos (nodes[243], nodes[558],  nodes[991]);
    nmos (nodes[493], nodes[1535],  nodes[859]);
    nmos (nodes[833], nodes[235],  nodes[859]);
    nmos (nodes[558], nodes[60],  nodes[1576]);
    nmos (nodes[558], nodes[84],  nodes[1576]);
    nmos (nodes[558], nodes[271],  nodes[1576]);
    nmos (nodes[558], nodes[370],  nodes[1576]);
    nmos (nodes[558], nodes[1612],  nodes[1576]);
    nmos (nodes[558], nodes[784],  nodes[1576]);
    nmos (nodes[558], nodes[204],  nodes[1576]);
    nmos (nodes[558], nodes[804],  nodes[1576]);
    nmos (nodes[558], nodes[1311],  nodes[1576]);
    nmos (nodes[558], nodes[1428],  nodes[1576]);
    nmos (nodes[558], nodes[492],  nodes[1576]);
    nmos (nodes[558], nodes[1204],  nodes[1576]);
    nmos (nodes[558], nodes[1259],  nodes[1576]);
    nmos (nodes[558], nodes[342],  nodes[1576]);
    nmos (nodes[558], nodes[857],  nodes[1576]);
    nmos (nodes[558], nodes[712],  nodes[1576]);
    nmos (nodes[558], nodes[776],  nodes[1576]);
    nmos (nodes[558], nodes[1168],  nodes[1576]);
    nmos (nodes[558], nodes[1721],  nodes[1576]);
    nmos (nodes[558], nodes[487],  nodes[1576]);
    nmos (nodes[558], nodes[579],  nodes[1576]);
    nmos (nodes[558], nodes[1239],  nodes[1576]);
    nmos (nodes[558], nodes[285],  nodes[1576]);
    nmos (nodes[558], nodes[1524],  nodes[1576]);
    nmos (nodes[558], nodes[0],  nodes[1576]);
    nmos (nodes[558], nodes[1478],  nodes[1576]);
    nmos (nodes[558], nodes[1210],  nodes[1576]);
    nmos (nodes[558], nodes[461],  nodes[1576]);
    nmos (nodes[558], nodes[660],  nodes[1576]);
    nmos (nodes[558], nodes[1557],  nodes[1576]);
    nmos (nodes[558], nodes[259],  nodes[1576]);
    nmos (nodes[558], nodes[352],  nodes[1576]);
    nmos (nodes[558], nodes[446],  nodes[1576]);
    nmos (nodes[558], nodes[528],  nodes[1576]);
    nmos (nodes[558], nodes[904],  nodes[1576]);
    nmos (nodes[558], nodes[1569],  nodes[1576]);
    nmos (nodes[558], nodes[1710],  nodes[1576]);
    nmos (nodes[558], nodes[219],  nodes[1576]);
    nmos (nodes[558], nodes[1385],  nodes[1576]);
    nmos (nodes[391], nodes[1147],  nodes[710]);
    nmos (nodes[991], nodes[1432],  nodes[859]);
    nmos (nodes[1302], nodes[96],  nodes[859]);
    nmos (nodes[704], nodes[1473],  nodes[859]);
    nmos (nodes[1503], nodes[1678],  nodes[859]);
    nmos (nodes[892], nodes[1645],  nodes[859]);
    nmos (nodes[558], nodes[806],  nodes[558]);
    nmos (nodes[578], nodes[589],  nodes[943]);
    nmos (nodes[558], nodes[1586],  nodes[682]);
    nmos (nodes[994], nodes[768],  nodes[943]);
    nmos (nodes[426], nodes[1386],  nodes[1316]);
    nmos (nodes[558], nodes[914],  nodes[1316]);
    nmos (nodes[413], nodes[657],  nodes[943]);
    nmos (nodes[780], nodes[1229],  nodes[943]);
    nmos (nodes[558], nodes[41],  nodes[1441]);
    nmos (nodes[1695], nodes[1318],  nodes[1535]);
    nmos (nodes[1398], nodes[558],  nodes[1535]);
    nmos (nodes[20], nodes[558],  nodes[1316]);
    nmos (nodes[387], nodes[558],  nodes[853]);
    nmos (nodes[558], nodes[670],  nodes[519]);
    nmos (nodes[670], nodes[558],  nodes[519]);
    nmos (nodes[1302], nodes[723],  nodes[283]);
    nmos (nodes[991], nodes[976],  nodes[283]);
    nmos (nodes[1647], nodes[493],  nodes[283]);
    nmos (nodes[1481], nodes[558],  nodes[698]);
    nmos (nodes[558], nodes[1371],  nodes[846]);
    nmos (nodes[558], nodes[333],  nodes[1201]);
    nmos (nodes[558], nodes[228],  nodes[21]);
    nmos (nodes[48], nodes[657],  nodes[21]);
    nmos (nodes[1110], nodes[1530],  nodes[943]);
    nmos (nodes[558], nodes[765],  nodes[1123]);
    nmos (nodes[558], nodes[661],  nodes[1607]);
    nmos (nodes[558], nodes[1178],  nodes[1652]);
    nmos (nodes[1225], nodes[1121],  nodes[943]);
    nmos (nodes[558], nodes[549],  nodes[1247]);
    nmos (nodes[558], nodes[783],  nodes[655]);
    nmos (nodes[558], nodes[227],  nodes[540]);
    nmos (nodes[558], nodes[1263],  nodes[602]);
    nmos (nodes[464], nodes[1661],  nodes[710]);
    nmos (nodes[558], nodes[255],  nodes[611]);
    nmos (nodes[657], nodes[741],  nodes[611]);
    nmos (nodes[558], nodes[917],  nodes[248]);
    nmos (nodes[513], nodes[558],  nodes[954]);
    nmos (nodes[322], nodes[558],  nodes[1026]);
    nmos (nodes[657], nodes[171],  nodes[1026]);
    nmos (nodes[1082], nodes[455],  nodes[1051]);
    nmos (nodes[1249], nodes[626],  nodes[1200]);
    nmos (nodes[191], nodes[456],  nodes[943]);
    nmos (nodes[1455], nodes[558],  nodes[822]);
    nmos (nodes[558], nodes[918],  nodes[404]);
    nmos (nodes[558], nodes[142],  nodes[404]);
    nmos (nodes[1331], nodes[558],  nodes[943]);
    nmos (nodes[1698], nodes[558],  nodes[943]);
    nmos (nodes[1479], nodes[558],  nodes[842]);
    nmos (nodes[66], nodes[657],  nodes[842]);
    nmos (nodes[1140], nodes[657],  nodes[713]);
    nmos (nodes[558], nodes[1231],  nodes[1409]);
    nmos (nodes[558], nodes[11],  nodes[1228]);
    nmos (nodes[558], nodes[1135],  nodes[166]);
    nmos (nodes[558], nodes[1695],  nodes[1522]);
    nmos (nodes[1398], nodes[558],  nodes[1522]);
    nmos (nodes[86], nodes[364],  nodes[943]);
    nmos (nodes[558], nodes[1117],  nodes[70]);
    nmos (nodes[558], nodes[10],  nodes[1211]);
    nmos (nodes[1308], nodes[558],  nodes[637]);
    nmos (nodes[657], nodes[349],  nodes[1608]);
    nmos (nodes[431], nodes[807],  nodes[1599]);
    nmos (nodes[1698], nodes[558],  nodes[1335]);
    nmos (nodes[558], nodes[252],  nodes[1665]);
    nmos (nodes[1263], nodes[558],  nodes[1247]);
    nmos (nodes[1489], nodes[1308],  nodes[1314]);
    nmos (nodes[558], nodes[637],  nodes[1314]);
    nmos (nodes[819], nodes[558],  nodes[596]);
    nmos (nodes[658], nodes[558],  nodes[565]);
    nmos (nodes[1383], nodes[1678],  nodes[1068]);
    nmos (nodes[351], nodes[235],  nodes[1068]);
    nmos (nodes[423], nodes[1535],  nodes[1068]);
    nmos (nodes[558], nodes[1294],  nodes[1605]);
    nmos (nodes[558], nodes[1112],  nodes[927]);
    nmos (nodes[558], nodes[1449],  nodes[958]);
    nmos (nodes[777], nodes[871],  nodes[943]);
    nmos (nodes[835], nodes[1229],  nodes[919]);
    nmos (nodes[1538], nodes[1486],  nodes[919]);
    nmos (nodes[200], nodes[558],  nodes[919]);
    nmos (nodes[558], nodes[1655],  nodes[1211]);
    nmos (nodes[809], nodes[558],  nodes[1077]);
    nmos (nodes[1410], nodes[558],  nodes[1077]);
    nmos (nodes[1668], nodes[705],  nodes[710]);
    nmos (nodes[558], nodes[1211],  nodes[273]);
    nmos (nodes[1445], nodes[558],  nodes[1492]);
    nmos (nodes[1457], nodes[558],  nodes[1492]);
    nmos (nodes[525], nodes[558],  nodes[266]);
    nmos (nodes[188], nodes[558],  nodes[1357]);
    nmos (nodes[123], nodes[246],  nodes[710]);
    nmos (nodes[657], nodes[7],  nodes[1415]);
    nmos (nodes[413], nodes[558],  nodes[217]);
    nmos (nodes[813], nodes[558],  nodes[440]);
    nmos (nodes[1280], nodes[558],  nodes[335]);
    nmos (nodes[558], nodes[1549],  nodes[1234]);
    nmos (nodes[558], nodes[851],  nodes[302]);
    nmos (nodes[94], nodes[1650],  nodes[710]);
    nmos (nodes[506], nodes[1602],  nodes[943]);
    nmos (nodes[853], nodes[558],  nodes[770]);
    nmos (nodes[558], nodes[163],  nodes[249]);
    nmos (nodes[558], nodes[1704],  nodes[249]);
    nmos (nodes[558], nodes[890],  nodes[1]);
    nmos (nodes[1601], nodes[558],  nodes[1329]);
    nmos (nodes[382], nodes[558],  nodes[1329]);
    nmos (nodes[1173], nodes[558],  nodes[1329]);
    nmos (nodes[1233], nodes[558],  nodes[1329]);
    nmos (nodes[1543], nodes[558],  nodes[1329]);
    nmos (nodes[76], nodes[558],  nodes[1329]);
    nmos (nodes[1540], nodes[558],  nodes[1329]);
    nmos (nodes[558], nodes[245],  nodes[1329]);
    nmos (nodes[786], nodes[558],  nodes[1329]);
    nmos (nodes[1482], nodes[558],  nodes[1329]);
    nmos (nodes[370], nodes[558],  nodes[1329]);
    nmos (nodes[552], nodes[558],  nodes[1329]);
    nmos (nodes[784], nodes[558],  nodes[1329]);
    nmos (nodes[1623], nodes[558],  nodes[1329]);
    nmos (nodes[403], nodes[558],  nodes[1329]);
    nmos (nodes[558], nodes[1311],  nodes[1329]);
    nmos (nodes[1355], nodes[558],  nodes[1329]);
    nmos (nodes[257], nodes[558],  nodes[1329]);
    nmos (nodes[179], nodes[558],  nodes[1329]);
    nmos (nodes[1086], nodes[558],  nodes[1329]);
    nmos (nodes[487], nodes[558],  nodes[1329]);
    nmos (nodes[145], nodes[558],  nodes[1329]);
    nmos (nodes[1478], nodes[558],  nodes[1329]);
    nmos (nodes[558], nodes[1557],  nodes[1329]);
    nmos (nodes[517], nodes[558],  nodes[1329]);
    nmos (nodes[352], nodes[558],  nodes[1329]);
    nmos (nodes[750], nodes[558],  nodes[1329]);
    nmos (nodes[932], nodes[558],  nodes[1329]);
    nmos (nodes[309], nodes[558],  nodes[1329]);
    nmos (nodes[1569], nodes[558],  nodes[1329]);
    nmos (nodes[301], nodes[558],  nodes[1329]);
    nmos (nodes[941], nodes[558],  nodes[199]);
    nmos (nodes[558], nodes[25],  nodes[256]);
    nmos (nodes[1059], nodes[633],  nodes[943]);
    nmos (nodes[40], nodes[1575],  nodes[943]);
    nmos (nodes[558], nodes[1554],  nodes[61]);
    nmos (nodes[479], nodes[558],  nodes[61]);
    nmos (nodes[558], nodes[485],  nodes[85]);
    nmos (nodes[558], nodes[679],  nodes[479]);
    nmos (nodes[558], nodes[1088],  nodes[873]);
    nmos (nodes[134], nodes[558],  nodes[259]);
    nmos (nodes[558], nodes[444],  nodes[823]);
    nmos (nodes[558], nodes[1433],  nodes[840]);
    nmos (nodes[381], nodes[657],  nodes[1315]);
    nmos (nodes[523], nodes[949],  nodes[83]);
    nmos (nodes[1406], nodes[558],  nodes[83]);
    nmos (nodes[558], nodes[570],  nodes[1220]);
    nmos (nodes[264], nodes[799],  nodes[943]);
    nmos (nodes[264], nodes[1693],  nodes[943]);
    nmos (nodes[558], nodes[46],  nodes[992]);
    nmos (nodes[252], nodes[558],  nodes[301]);
    nmos (nodes[241], nodes[558],  nodes[745]);
    nmos (nodes[1446], nodes[558],  nodes[771]);
    nmos (nodes[465], nodes[430],  nodes[771]);
    nmos (nodes[766], nodes[474],  nodes[1184]);
    nmos (nodes[410], nodes[558],  nodes[1184]);
    nmos (nodes[558], nodes[1671],  nodes[1077]);
    nmos (nodes[1460], nodes[558],  nodes[1077]);
    nmos (nodes[558], nodes[811],  nodes[838]);
    nmos (nodes[26], nodes[558],  nodes[1112]);
    nmos (nodes[209], nodes[558],  nodes[113]);
    nmos (nodes[759], nodes[187],  nodes[710]);
    nmos (nodes[558], nodes[1687],  nodes[1108]);
    nmos (nodes[1035], nodes[558],  nodes[943]);
    nmos (nodes[1328], nodes[558],  nodes[541]);
    nmos (nodes[1150], nodes[872],  nodes[129]);
    nmos (nodes[558], nodes[587],  nodes[1283]);
    nmos (nodes[54], nodes[401],  nodes[129]);
    nmos (nodes[1109], nodes[558],  nodes[902]);
    nmos (nodes[1109], nodes[558],  nodes[902]);
    nmos (nodes[1289], nodes[558],  nodes[902]);
    nmos (nodes[558], nodes[1047],  nodes[830]);
    nmos (nodes[657], nodes[534],  nodes[830]);
    nmos (nodes[766], nodes[558],  nodes[1643]);
    nmos (nodes[558], nodes[1704],  nodes[1643]);
    nmos (nodes[410], nodes[558],  nodes[1643]);
    nmos (nodes[1587], nodes[558],  nodes[1077]);
    nmos (nodes[540], nodes[558],  nodes[1077]);
    nmos (nodes[1000], nodes[1408],  nodes[1044]);
    nmos (nodes[215], nodes[1379],  nodes[943]);
    nmos (nodes[345], nodes[1279],  nodes[986]);
    nmos (nodes[1108], nodes[1722],  nodes[247]);
    nmos (nodes[209], nodes[991],  nodes[247]);
    nmos (nodes[1496], nodes[1473],  nodes[247]);
    nmos (nodes[1302], nodes[141],  nodes[247]);
    nmos (nodes[892], nodes[27],  nodes[247]);
    nmos (nodes[1503], nodes[1301],  nodes[247]);
    nmos (nodes[652], nodes[833],  nodes[247]);
    nmos (nodes[1206], nodes[493],  nodes[247]);
    nmos (nodes[869], nodes[1128],  nodes[943]);
    nmos (nodes[558], nodes[772],  nodes[1674]);
    nmos (nodes[558], nodes[446],  nodes[909]);
    nmos (nodes[558], nodes[528],  nodes[909]);
    nmos (nodes[558], nodes[0],  nodes[909]);
    nmos (nodes[558], nodes[1210],  nodes[909]);
    nmos (nodes[558], nodes[1385],  nodes[909]);
    nmos (nodes[558], nodes[370],  nodes[909]);
    nmos (nodes[558], nodes[784],  nodes[909]);
    nmos (nodes[558], nodes[776],  nodes[909]);
    nmos (nodes[558], nodes[1168],  nodes[909]);
    nmos (nodes[1221], nodes[104],  nodes[943]);
    nmos (nodes[1186], nodes[558],  nodes[943]);
    nmos (nodes[558], nodes[1263],  nodes[943]);
    nmos (nodes[325], nodes[558],  nodes[943]);
    nmos (nodes[801], nodes[558],  nodes[943]);
    nmos (nodes[420], nodes[47],  nodes[710]);
    nmos (nodes[1706], nodes[558],  nodes[937]);
    nmos (nodes[1704], nodes[558],  nodes[937]);
    nmos (nodes[1345], nodes[558],  nodes[937]);
    nmos (nodes[558], nodes[717],  nodes[1132]);
    nmos (nodes[1380], nodes[666],  nodes[710]);
    nmos (nodes[558], nodes[334],  nodes[1382]);
    nmos (nodes[657], nodes[676],  nodes[617]);
    nmos (nodes[527], nodes[1474],  nodes[710]);
    nmos (nodes[558], nodes[1705],  nodes[630]);
    nmos (nodes[558], nodes[898],  nodes[1518]);
    nmos (nodes[558], nodes[1710],  nodes[996]);
    nmos (nodes[1601], nodes[558],  nodes[996]);
    nmos (nodes[382], nodes[558],  nodes[996]);
    nmos (nodes[1173], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[1233],  nodes[996]);
    nmos (nodes[558], nodes[1658],  nodes[996]);
    nmos (nodes[558], nodes[1664],  nodes[996]);
    nmos (nodes[558], nodes[1482],  nodes[996]);
    nmos (nodes[558], nodes[665],  nodes[996]);
    nmos (nodes[286], nodes[558],  nodes[996]);
    nmos (nodes[271], nodes[558],  nodes[996]);
    nmos (nodes[370], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[552],  nodes[996]);
    nmos (nodes[558], nodes[1612],  nodes[996]);
    nmos (nodes[558], nodes[1487],  nodes[996]);
    nmos (nodes[558], nodes[784],  nodes[996]);
    nmos (nodes[558], nodes[764],  nodes[996]);
    nmos (nodes[1582], nodes[558],  nodes[996]);
    nmos (nodes[1031], nodes[558],  nodes[996]);
    nmos (nodes[804], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[1311],  nodes[996]);
    nmos (nodes[558], nodes[1520],  nodes[996]);
    nmos (nodes[558], nodes[857],  nodes[996]);
    nmos (nodes[558], nodes[712],  nodes[996]);
    nmos (nodes[558], nodes[1337],  nodes[996]);
    nmos (nodes[1381], nodes[558],  nodes[996]);
    nmos (nodes[776], nodes[558],  nodes[996]);
    nmos (nodes[157], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[257],  nodes[996]);
    nmos (nodes[558], nodes[131],  nodes[996]);
    nmos (nodes[558], nodes[4],  nodes[996]);
    nmos (nodes[558], nodes[303],  nodes[996]);
    nmos (nodes[558], nodes[1721],  nodes[996]);
    nmos (nodes[1086], nodes[558],  nodes[996]);
    nmos (nodes[487], nodes[558],  nodes[996]);
    nmos (nodes[579], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[1239],  nodes[996]);
    nmos (nodes[558], nodes[0],  nodes[996]);
    nmos (nodes[558], nodes[1478],  nodes[996]);
    nmos (nodes[558], nodes[594],  nodes[996]);
    nmos (nodes[558], nodes[660],  nodes[996]);
    nmos (nodes[1557], nodes[558],  nodes[996]);
    nmos (nodes[259], nodes[558],  nodes[996]);
    nmos (nodes[1052], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[791],  nodes[996]);
    nmos (nodes[558], nodes[352],  nodes[996]);
    nmos (nodes[558], nodes[750],  nodes[996]);
    nmos (nodes[558], nodes[932],  nodes[996]);
    nmos (nodes[558], nodes[1589],  nodes[996]);
    nmos (nodes[446], nodes[558],  nodes[996]);
    nmos (nodes[528], nodes[558],  nodes[996]);
    nmos (nodes[309], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[1430],  nodes[996]);
    nmos (nodes[558], nodes[1292],  nodes[996]);
    nmos (nodes[558], nodes[1646],  nodes[996]);
    nmos (nodes[558], nodes[1114],  nodes[996]);
    nmos (nodes[558], nodes[1476],  nodes[996]);
    nmos (nodes[1226], nodes[558],  nodes[996]);
    nmos (nodes[1569], nodes[558],  nodes[996]);
    nmos (nodes[950], nodes[558],  nodes[996]);
    nmos (nodes[558], nodes[1050],  nodes[996]);
    nmos (nodes[558], nodes[1419],  nodes[996]);
    nmos (nodes[558], nodes[1164],  nodes[996]);
    nmos (nodes[558], nodes[995],  nodes[312]);
    nmos (nodes[742], nodes[854],  nodes[312]);
    nmos (nodes[558], nodes[1425],  nodes[988]);
    nmos (nodes[1382], nodes[1291],  nodes[710]);
    nmos (nodes[926], nodes[558],  nodes[717]);
    nmos (nodes[1087], nodes[558],  nodes[717]);
    nmos (nodes[1545], nodes[558],  nodes[1034]);
    nmos (nodes[657], nodes[994],  nodes[1034]);
    nmos (nodes[1410], nodes[558],  nodes[1690]);
    nmos (nodes[744], nodes[558],  nodes[1302]);
    nmos (nodes[558], nodes[1558],  nodes[40]);
    nmos (nodes[12], nodes[558],  nodes[40]);
    nmos (nodes[1016], nodes[558],  nodes[1282]);
    nmos (nodes[558], nodes[551],  nodes[393]);
    nmos (nodes[1085], nodes[596],  nodes[943]);
    nmos (nodes[685], nodes[1175],  nodes[943]);
    nmos (nodes[558], nodes[1312],  nodes[1291]);
    nmos (nodes[532], nodes[1013],  nodes[592]);
    nmos (nodes[1217], nodes[558],  nodes[592]);
    nmos (nodes[558], nodes[1510],  nodes[1021]);
    nmos (nodes[558], nodes[365],  nodes[809]);
    nmos (nodes[77], nodes[558],  nodes[90]);
    nmos (nodes[558], nodes[1454],  nodes[852]);
    nmos (nodes[558], nodes[260],  nodes[852]);
    nmos (nodes[1555], nodes[1107],  nodes[324]);
    nmos (nodes[1325], nodes[558],  nodes[769]);
    nmos (nodes[1072], nodes[657],  nodes[769]);
    nmos (nodes[1643], nodes[558],  nodes[900]);
    nmos (nodes[1393], nodes[1393],  nodes[147]);
    nmos (nodes[558], nodes[1393],  nodes[147]);
    nmos (nodes[558], nodes[1393],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[1393], nodes[558],  nodes[147]);
    nmos (nodes[558], nodes[1376],  nodes[1473]);
    nmos (nodes[125], nodes[558],  nodes[365]);
    nmos (nodes[558], nodes[363],  nodes[537]);
    nmos (nodes[558], nodes[731],  nodes[993]);
    nmos (nodes[1203], nodes[263],  nodes[753]);
    nmos (nodes[1629], nodes[558],  nodes[753]);
    nmos (nodes[558], nodes[827],  nodes[926]);
    nmos (nodes[339], nodes[632],  nodes[943]);
    nmos (nodes[108], nodes[558],  nodes[1364]);
    nmos (nodes[1666], nodes[657],  nodes[1364]);
    nmos (nodes[953], nodes[558],  nodes[425]);
    nmos (nodes[558], nodes[943],  nodes[1467]);
    nmos (nodes[558], nodes[943],  nodes[1467]);
    nmos (nodes[558], nodes[943],  nodes[1467]);
    nmos (nodes[943], nodes[558],  nodes[1467]);
    nmos (nodes[720], nodes[558],  nodes[56]);
    nmos (nodes[1494], nodes[558],  nodes[260]);
    nmos (nodes[558], nodes[1009],  nodes[735]);
    nmos (nodes[558], nodes[935],  nodes[1242]);
    nmos (nodes[146], nodes[558],  nodes[5]);
    nmos (nodes[558], nodes[438],  nodes[1462]);
    nmos (nodes[558], nodes[1544],  nodes[1115]);
    nmos (nodes[1658], nodes[558],  nodes[1394]);
    nmos (nodes[985], nodes[558],  nodes[1394]);
    nmos (nodes[1664], nodes[558],  nodes[1394]);
    nmos (nodes[682], nodes[558],  nodes[1394]);
    nmos (nodes[665], nodes[558],  nodes[1394]);
    nmos (nodes[286], nodes[558],  nodes[1394]);
    nmos (nodes[271], nodes[558],  nodes[1394]);
    nmos (nodes[1612], nodes[558],  nodes[1394]);
    nmos (nodes[1487], nodes[558],  nodes[1394]);
    nmos (nodes[244], nodes[558],  nodes[1394]);
    nmos (nodes[1520], nodes[558],  nodes[1394]);
    nmos (nodes[324], nodes[558],  nodes[1394]);
    nmos (nodes[712], nodes[558],  nodes[1394]);
    nmos (nodes[787], nodes[558],  nodes[1394]);
    nmos (nodes[575], nodes[558],  nodes[1394]);
    nmos (nodes[1466], nodes[558],  nodes[1394]);
    nmos (nodes[776], nodes[558],  nodes[1394]);
    nmos (nodes[822], nodes[558],  nodes[1394]);
    nmos (nodes[131], nodes[558],  nodes[1394]);
    nmos (nodes[1420], nodes[558],  nodes[1394]);
    nmos (nodes[4], nodes[558],  nodes[1394]);
    nmos (nodes[167], nodes[558],  nodes[1394]);
    nmos (nodes[303], nodes[558],  nodes[1394]);
    nmos (nodes[1504], nodes[558],  nodes[1394]);
    nmos (nodes[579], nodes[558],  nodes[1394]);
    nmos (nodes[0], nodes[558],  nodes[1394]);
    nmos (nodes[259], nodes[558],  nodes[1394]);
    nmos (nodes[528], nodes[558],  nodes[1394]);
    nmos (nodes[1430], nodes[558],  nodes[1394]);
    nmos (nodes[1646], nodes[558],  nodes[1394]);
    nmos (nodes[1155], nodes[558],  nodes[1394]);
    nmos (nodes[1476], nodes[558],  nodes[1394]);
    nmos (nodes[1226], nodes[558],  nodes[1394]);
    nmos (nodes[1164], nodes[558],  nodes[1394]);
    nmos (nodes[558], nodes[1497],  nodes[1438]);
    nmos (nodes[558], nodes[887],  nodes[1254]);
    nmos (nodes[887], nodes[558],  nodes[1254]);
    nmos (nodes[887], nodes[558],  nodes[1254]);
    nmos (nodes[887], nodes[558],  nodes[1254]);
    nmos (nodes[558], nodes[302],  nodes[540]);
    nmos (nodes[365], nodes[558],  nodes[540]);
    nmos (nodes[558], nodes[1294],  nodes[540]);
    nmos (nodes[506], nodes[558],  nodes[236]);
    nmos (nodes[558], nodes[1656],  nodes[1580]);
    nmos (nodes[558], nodes[1159],  nodes[1580]);
    nmos (nodes[1550], nodes[845],  nodes[1573]);
    nmos (nodes[558], nodes[959],  nodes[430]);
    nmos (nodes[166], nodes[578],  nodes[1263]);
    nmos (nodes[1336], nodes[1724],  nodes[1263]);
    nmos (nodes[574], nodes[558],  nodes[1256]);
    nmos (nodes[1287], nodes[1694],  nodes[1263]);
    nmos (nodes[1188], nodes[242],  nodes[1263]);
    nmos (nodes[1405], nodes[436],  nodes[1263]);
    nmos (nodes[520], nodes[558],  nodes[224]);
    nmos (nodes[37], nodes[657],  nodes[224]);
    nmos (nodes[831], nodes[558],  nodes[1719]);
    nmos (nodes[570], nodes[558],  nodes[1144]);
    nmos (nodes[558], nodes[1394],  nodes[1329]);
    nmos (nodes[879], nodes[558],  nodes[248]);
    nmos (nodes[538], nodes[558],  nodes[1599]);
    nmos (nodes[399], nodes[657],  nodes[1296]);
    nmos (nodes[1599], nodes[558],  nodes[103]);
    nmos (nodes[1577], nodes[1391],  nodes[943]);
    nmos (nodes[1255], nodes[558],  nodes[531]);
    nmos (nodes[59], nodes[657],  nodes[531]);
    nmos (nodes[298], nodes[657],  nodes[63]);
    nmos (nodes[999], nodes[668],  nodes[943]);
    nmos (nodes[907], nodes[1298],  nodes[821]);
    nmos (nodes[1404], nodes[1106],  nodes[943]);
    nmos (nodes[240], nodes[558],  nodes[498]);
    nmos (nodes[240], nodes[558],  nodes[498]);
    nmos (nodes[240], nodes[558],  nodes[498]);
    nmos (nodes[1464], nodes[558],  nodes[1612]);
    nmos (nodes[1649], nodes[558],  nodes[712]);
    nmos (nodes[1150], nodes[767],  nodes[801]);
    nmos (nodes[189], nodes[841],  nodes[1432]);
    nmos (nodes[155], nodes[558],  nodes[1432]);
    nmos (nodes[558], nodes[1186],  nodes[662]);
    nmos (nodes[33], nodes[558],  nodes[469]);
    nmos (nodes[558], nodes[86],  nodes[1232]);
    nmos (nodes[1676], nodes[558],  nodes[1232]);
    nmos (nodes[657], nodes[634],  nodes[1232]);
    nmos (nodes[1709], nodes[558],  nodes[1434]);
    nmos (nodes[1389], nodes[558],  nodes[752]);
    nmos (nodes[216], nodes[558],  nodes[681]);
    nmos (nodes[558], nodes[639],  nodes[130]);
    nmos (nodes[558], nodes[104],  nodes[275]);
    nmos (nodes[851], nodes[1515],  nodes[1019]);
    nmos (nodes[558], nodes[231],  nodes[1019]);
    nmos (nodes[558], nodes[1458],  nodes[731]);
    nmos (nodes[1120], nodes[558],  nodes[248]);
    nmos (nodes[2], nodes[1039],  nodes[248]);
    nmos (nodes[300], nodes[558],  nodes[342]);
    nmos (nodes[558], nodes[117],  nodes[1398]);
    nmos (nodes[1241], nodes[558],  nodes[1398]);
    nmos (nodes[1140], nodes[558],  nodes[617]);
    nmos (nodes[558], nodes[1295],  nodes[1527]);
    nmos (nodes[558], nodes[1515],  nodes[125]);
    nmos (nodes[90], nodes[558],  nodes[1625]);
    nmos (nodes[558], nodes[1379],  nodes[1476]);
    nmos (nodes[558], nodes[275],  nodes[1697]);
    nmos (nodes[595], nodes[558],  nodes[1168]);
    nmos (nodes[558], nodes[623],  nodes[143]);
    nmos (nodes[558], nodes[1347],  nodes[782]);
    nmos (nodes[558], nodes[934],  nodes[366]);
    nmos (nodes[72], nodes[622],  nodes[898]);
    nmos (nodes[208], nodes[900],  nodes[898]);
    nmos (nodes[1647], nodes[1611],  nodes[898]);
    nmos (nodes[1458], nodes[377],  nodes[898]);
    nmos (nodes[976], nodes[1022],  nodes[898]);
    nmos (nodes[488], nodes[1139],  nodes[898]);
    nmos (nodes[723], nodes[1359],  nodes[898]);
    nmos (nodes[481], nodes[655],  nodes[898]);
    nmos (nodes[166], nodes[483],  nodes[140]);
    nmos (nodes[121], nodes[618],  nodes[1468]);
    nmos (nodes[254], nodes[558],  nodes[483]);
    nmos (nodes[1038], nodes[558],  nodes[336]);
    nmos (nodes[1158], nodes[515],  nodes[1542]);
    nmos (nodes[1253], nodes[558],  nodes[1542]);
    nmos (nodes[558], nodes[984],  nodes[1247]);
    nmos (nodes[870], nodes[558],  nodes[576]);
    nmos (nodes[870], nodes[558],  nodes[576]);
    nmos (nodes[870], nodes[558],  nodes[576]);
    nmos (nodes[515], nodes[558],  nodes[1253]);
    nmos (nodes[160], nodes[558],  nodes[934]);
    nmos (nodes[558], nodes[1689],  nodes[837]);
    nmos (nodes[910], nodes[558],  nodes[590]);
    nmos (nodes[54], nodes[332],  nodes[1700]);
    nmos (nodes[423], nodes[558],  nodes[493]);
    nmos (nodes[774], nodes[974],  nodes[943]);
    nmos (nodes[968], nodes[934],  nodes[943]);
    nmos (nodes[415], nodes[1196],  nodes[943]);
    nmos (nodes[1688], nodes[680],  nodes[943]);
    nmos (nodes[558], nodes[106],  nodes[1528]);
    nmos (nodes[669], nodes[558],  nodes[303]);
    nmos (nodes[235], nodes[121],  nodes[437]);
    nmos (nodes[1535], nodes[1299],  nodes[437]);
    nmos (nodes[657], nodes[349],  nodes[1608]);
    nmos (nodes[1432], nodes[1282],  nodes[437]);
    nmos (nodes[1645], nodes[1437],  nodes[437]);
    nmos (nodes[1630], nodes[1678],  nodes[437]);
    nmos (nodes[1465], nodes[1126],  nodes[943]);
    nmos (nodes[96], nodes[684],  nodes[437]);
    nmos (nodes[899], nodes[19],  nodes[943]);
    nmos (nodes[1179], nodes[558],  nodes[725]);
    nmos (nodes[558], nodes[1286],  nodes[930]);
    nmos (nodes[718], nodes[558],  nodes[1005]);
    nmos (nodes[558], nodes[1591],  nodes[558]);
    nmos (nodes[978], nodes[1618],  nodes[943]);
    nmos (nodes[111], nodes[558],  nodes[945]);
    nmos (nodes[1123], nodes[304],  nodes[943]);
    nmos (nodes[558], nodes[896],  nodes[650]);
    nmos (nodes[558], nodes[1211],  nodes[1002]);
    nmos (nodes[299], nodes[1470],  nodes[1416]);
    nmos (nodes[558], nodes[152],  nodes[952]);
    nmos (nodes[272], nodes[558],  nodes[862]);
    nmos (nodes[1351], nodes[1717],  nodes[258]);
    nmos (nodes[1150], nodes[1709],  nodes[1263]);
    nmos (nodes[558], nodes[1228],  nodes[669]);
    nmos (nodes[558], nodes[1393],  nodes[558]);
    nmos (nodes[1252], nodes[1374],  nodes[943]);
    nmos (nodes[558], nodes[1483],  nodes[1627]);
    nmos (nodes[1084], nodes[558],  nodes[1627]);
    nmos (nodes[558], nodes[1707],  nodes[936]);
    nmos (nodes[558], nodes[388],  nodes[936]);
    nmos (nodes[1344], nodes[727],  nodes[943]);
    nmos (nodes[1265], nodes[558],  nodes[502]);
    nmos (nodes[1251], nodes[558],  nodes[1640]);
    nmos (nodes[420], nodes[558],  nodes[865]);
    nmos (nodes[558], nodes[645],  nodes[1032]);
    nmos (nodes[558], nodes[60],  nodes[1384]);
    nmos (nodes[558], nodes[1512],  nodes[1384]);
    nmos (nodes[558], nodes[382],  nodes[1384]);
    nmos (nodes[558], nodes[1173],  nodes[1384]);
    nmos (nodes[558], nodes[84],  nodes[1384]);
    nmos (nodes[558], nodes[1543],  nodes[1384]);
    nmos (nodes[558], nodes[76],  nodes[1384]);
    nmos (nodes[558], nodes[245],  nodes[1384]);
    nmos (nodes[558], nodes[786],  nodes[1384]);
    nmos (nodes[558], nodes[1664],  nodes[1384]);
    nmos (nodes[558], nodes[682],  nodes[1384]);
    nmos (nodes[558], nodes[1482],  nodes[1384]);
    nmos (nodes[558], nodes[271],  nodes[1384]);
    nmos (nodes[558], nodes[370],  nodes[1384]);
    nmos (nodes[558], nodes[552],  nodes[1384]);
    nmos (nodes[558], nodes[1612],  nodes[1384]);
    nmos (nodes[558], nodes[1487],  nodes[1384]);
    nmos (nodes[558], nodes[784],  nodes[1384]);
    nmos (nodes[558], nodes[1582],  nodes[1384]);
    nmos (nodes[558], nodes[804],  nodes[1384]);
    nmos (nodes[558], nodes[1311],  nodes[1384]);
    nmos (nodes[558], nodes[1428],  nodes[1384]);
    nmos (nodes[558], nodes[492],  nodes[1384]);
    nmos (nodes[558], nodes[1204],  nodes[1384]);
    nmos (nodes[558], nodes[1520],  nodes[1384]);
    nmos (nodes[558], nodes[1259],  nodes[1384]);
    nmos (nodes[558], nodes[342],  nodes[1384]);
    nmos (nodes[558], nodes[857],  nodes[1384]);
    nmos (nodes[558], nodes[712],  nodes[1384]);
    nmos (nodes[558], nodes[776],  nodes[1384]);
    nmos (nodes[558], nodes[157],  nodes[1384]);
    nmos (nodes[558], nodes[257],  nodes[1384]);
    nmos (nodes[558], nodes[1324],  nodes[1384]);
    nmos (nodes[558], nodes[179],  nodes[1384]);
    nmos (nodes[558], nodes[131],  nodes[1384]);
    nmos (nodes[558], nodes[4],  nodes[1384]);
    nmos (nodes[558], nodes[1396],  nodes[1384]);
    nmos (nodes[558], nodes[167],  nodes[1384]);
    nmos (nodes[558], nodes[1168],  nodes[1384]);
    nmos (nodes[558], nodes[1721],  nodes[1384]);
    nmos (nodes[558], nodes[1086],  nodes[1384]);
    nmos (nodes[558], nodes[1074],  nodes[1384]);
    nmos (nodes[558], nodes[487],  nodes[1384]);
    nmos (nodes[558], nodes[579],  nodes[1384]);
    nmos (nodes[558], nodes[1239],  nodes[1384]);
    nmos (nodes[558], nodes[1524],  nodes[1384]);
    nmos (nodes[558], nodes[0],  nodes[1384]);
    nmos (nodes[558], nodes[1478],  nodes[1384]);
    nmos (nodes[558], nodes[1210],  nodes[1384]);
    nmos (nodes[558], nodes[461],  nodes[1384]);
    nmos (nodes[558], nodes[660],  nodes[1384]);
    nmos (nodes[558], nodes[1557],  nodes[1384]);
    nmos (nodes[558], nodes[259],  nodes[1384]);
    nmos (nodes[558], nodes[791],  nodes[1384]);
    nmos (nodes[558], nodes[352],  nodes[1384]);
    nmos (nodes[558], nodes[750],  nodes[1384]);
    nmos (nodes[558], nodes[932],  nodes[1384]);
    nmos (nodes[558], nodes[446],  nodes[1384]);
    nmos (nodes[558], nodes[528],  nodes[1384]);
    nmos (nodes[558], nodes[1430],  nodes[1384]);
    nmos (nodes[558], nodes[1292],  nodes[1384]);
    nmos (nodes[558], nodes[1114],  nodes[1384]);
    nmos (nodes[558], nodes[1226],  nodes[1384]);
    nmos (nodes[558], nodes[1569],  nodes[1384]);
    nmos (nodes[558], nodes[1665],  nodes[1384]);
    nmos (nodes[558], nodes[1050],  nodes[1384]);
    nmos (nodes[558], nodes[1419],  nodes[1384]);
    nmos (nodes[558], nodes[1385],  nodes[1384]);
    nmos (nodes[558], nodes[1164],  nodes[1384]);
    nmos (nodes[558], nodes[1006],  nodes[1384]);
    nmos (nodes[45], nodes[1712],  nodes[943]);
    nmos (nodes[871], nodes[558],  nodes[1561]);
    nmos (nodes[558], nodes[726],  nodes[1210]);
    nmos (nodes[256], nodes[558],  nodes[1210]);
    nmos (nodes[1076], nodes[558],  nodes[1463]);
    nmos (nodes[147], nodes[657],  nodes[1463]);
    nmos (nodes[1711], nodes[558],  nodes[183]);
    nmos (nodes[1455], nodes[558],  nodes[257]);
    nmos (nodes[564], nodes[64],  nodes[943]);
    nmos (nodes[429], nodes[659],  nodes[943]);
    nmos (nodes[558], nodes[1209],  nodes[1213]);
    nmos (nodes[48], nodes[558],  nodes[228]);
    nmos (nodes[186], nodes[558],  nodes[1224]);
    nmos (nodes[1414], nodes[558],  nodes[495]);
    nmos (nodes[1441], nodes[558],  nodes[1277]);
    nmos (nodes[41], nodes[657],  nodes[1277]);
    nmos (nodes[781], nodes[558],  nodes[248]);
    nmos (nodes[781], nodes[558],  nodes[248]);
    nmos (nodes[558], nodes[930],  nodes[134]);
    nmos (nodes[558], nodes[467],  nodes[134]);
    nmos (nodes[67], nodes[449],  nodes[943]);
    nmos (nodes[558], nodes[1080],  nodes[811]);
    nmos (nodes[100], nodes[1205],  nodes[811]);
    nmos (nodes[657], nodes[991],  nodes[943]);
    nmos (nodes[1641], nodes[558],  nodes[809]);
    nmos (nodes[1547], nodes[1192],  nodes[609]);
    nmos (nodes[1264], nodes[1209],  nodes[609]);
    nmos (nodes[384], nodes[558],  nodes[1412]);
    nmos (nodes[558], nodes[62],  nodes[1349]);
    nmos (nodes[720], nodes[1338],  nodes[710]);
    nmos (nodes[1109], nodes[558],  nodes[1464]);
    nmos (nodes[703], nodes[227],  nodes[710]);
    nmos (nodes[657], nodes[166],  nodes[943]);
    nmos (nodes[181], nodes[548],  nodes[943]);
    nmos (nodes[1306], nodes[1095],  nodes[710]);
    nmos (nodes[43], nodes[558],  nodes[710]);
    nmos (nodes[839], nodes[558],  nodes[710]);
    nmos (nodes[507], nodes[558],  nodes[1049]);
    nmos (nodes[954], nodes[558],  nodes[338]);
    nmos (nodes[1522], nodes[1001],  nodes[549]);
    nmos (nodes[558], nodes[981],  nodes[615]);
    nmos (nodes[558], nodes[1260],  nodes[598]);
    nmos (nodes[328], nodes[558],  nodes[310]);
    nmos (nodes[558], nodes[494],  nodes[1539]);
    nmos (nodes[657], nodes[13],  nodes[943]);
    nmos (nodes[1299], nodes[657],  nodes[943]);
    nmos (nodes[558], nodes[501],  nodes[180]);
    nmos (nodes[558], nodes[976],  nodes[1102]);
    nmos (nodes[192], nodes[239],  nodes[1048]);
    nmos (nodes[1531], nodes[558],  nodes[184]);
    nmos (nodes[1485], nodes[1199],  nodes[943]);
    nmos (nodes[56], nodes[824],  nodes[943]);
    nmos (nodes[558], nodes[886],  nodes[943]);
    nmos (nodes[1307], nodes[524],  nodes[639]);
    nmos (nodes[28], nodes[577],  nodes[639]);
    nmos (nodes[364], nodes[738],  nodes[639]);
    nmos (nodes[1513], nodes[463],  nodes[639]);
    nmos (nodes[558], nodes[1094],  nodes[1630]);
    nmos (nodes[1712], nodes[558],  nodes[264]);
    nmos (nodes[558], nodes[261],  nodes[461]);
    nmos (nodes[558], nodes[726],  nodes[461]);
    nmos (nodes[1077], nodes[380],  nodes[879]);
    nmos (nodes[558], nodes[238],  nodes[1713]);
    nmos (nodes[1354], nodes[623],  nodes[1628]);
    nmos (nodes[713], nodes[558],  nodes[907]);
    nmos (nodes[1282], nodes[1022],  nodes[414]);
    nmos (nodes[1139], nodes[413],  nodes[414]);
    nmos (nodes[684], nodes[1359],  nodes[414]);
    nmos (nodes[655], nodes[1242],  nodes[414]);
    nmos (nodes[1630], nodes[622],  nodes[414]);
    nmos (nodes[900], nodes[1437],  nodes[414]);
    nmos (nodes[377], nodes[121],  nodes[414]);
    nmos (nodes[1185], nodes[558],  nodes[248]);
    nmos (nodes[744], nodes[558],  nodes[1108]);
    nmos (nodes[558], nodes[140],  nodes[1271]);
    nmos (nodes[312], nodes[558],  nodes[159]);
    nmos (nodes[1287], nodes[1637],  nodes[129]);
    nmos (nodes[1659], nodes[558],  nodes[499]);
    nmos (nodes[743], nodes[558],  nodes[499]);
    nmos (nodes[558], nodes[252],  nodes[950]);
    nmos (nodes[618], nodes[558],  nodes[1029]);
    nmos (nodes[695], nodes[1341],  nodes[943]);
    nmos (nodes[657], nodes[1237],  nodes[475]);
    nmos (nodes[1001], nodes[1435],  nodes[874]);
    nmos (nodes[558], nodes[1340],  nodes[642]);
    nmos (nodes[558], nodes[1340],  nodes[642]);
    nmos (nodes[558], nodes[1340],  nodes[642]);
    nmos (nodes[558], nodes[1340],  nodes[642]);
    nmos (nodes[558], nodes[152],  nodes[1002]);
    nmos (nodes[1407], nodes[558],  nodes[572]);
    nmos (nodes[334], nodes[1078],  nodes[943]);
    nmos (nodes[657], nodes[451],  nodes[1479]);
    nmos (nodes[657], nodes[451],  nodes[1479]);
    nmos (nodes[657], nodes[451],  nodes[1479]);
    nmos (nodes[451], nodes[657],  nodes[1479]);
    nmos (nodes[657], nodes[451],  nodes[1479]);
    nmos (nodes[1521], nodes[558],  nodes[1648]);
    nmos (nodes[558], nodes[14],  nodes[323]);
    nmos (nodes[593], nodes[558],  nodes[355]);
    nmos (nodes[1700], nodes[657],  nodes[355]);
    nmos (nodes[558], nodes[814],  nodes[392]);
    nmos (nodes[558], nodes[557],  nodes[392]);
    nmos (nodes[558], nodes[82],  nodes[794]);
    nmos (nodes[558], nodes[82],  nodes[794]);
    nmos (nodes[82], nodes[558],  nodes[794]);
    nmos (nodes[82], nodes[558],  nodes[794]);
    nmos (nodes[558], nodes[82],  nodes[794]);
    nmos (nodes[558], nodes[82],  nodes[794]);
    nmos (nodes[558], nodes[82],  nodes[794]);
    nmos (nodes[1436], nodes[1155],  nodes[943]);
    nmos (nodes[610], nodes[696],  nodes[943]);
    nmos (nodes[558], nodes[811],  nodes[1146]);
    nmos (nodes[558], nodes[1440],  nodes[248]);
    nmos (nodes[936], nodes[558],  nodes[841]);
    nmos (nodes[558], nodes[1501],  nodes[63]);
    nmos (nodes[558], nodes[23],  nodes[63]);
    nmos (nodes[558], nodes[801],  nodes[1247]);
    nmos (nodes[558], nodes[1230],  nodes[43]);
    nmos (nodes[558], nodes[570],  nodes[122]);
    nmos (nodes[558], nodes[1313],  nodes[649]);
    nmos (nodes[558], nodes[640],  nodes[649]);
    nmos (nodes[558], nodes[452],  nodes[1332]);
    nmos (nodes[558], nodes[1691],  nodes[1332]);
    nmos (nodes[558], nodes[1196],  nodes[934]);
    nmos (nodes[1585], nodes[558],  nodes[943]);
    nmos (nodes[1518], nodes[558],  nodes[1270]);
    nmos (nodes[657], nodes[898],  nodes[1270]);
    nmos (nodes[558], nodes[432],  nodes[1188]);
    nmos (nodes[558], nodes[432],  nodes[1188]);
    nmos (nodes[714], nodes[558],  nodes[906]);
    nmos (nodes[214], nodes[558],  nodes[906]);
    nmos (nodes[578], nodes[558],  nodes[1017]);
    nmos (nodes[558], nodes[462],  nodes[1338]);
    nmos (nodes[558], nodes[1350],  nodes[1382]);
    nmos (nodes[1591], nodes[657],  nodes[7]);
    nmos (nodes[1591], nodes[657],  nodes[7]);
    nmos (nodes[1591], nodes[657],  nodes[7]);
    nmos (nodes[1526], nodes[558],  nodes[680]);
    nmos (nodes[760], nodes[629],  nodes[943]);
    nmos (nodes[1427], nodes[558],  nodes[967]);
    nmos (nodes[558], nodes[852],  nodes[1001]);
    nmos (nodes[558], nodes[852],  nodes[1001]);
    nmos (nodes[558], nodes[211],  nodes[138]);
    nmos (nodes[558], nodes[211],  nodes[138]);
    nmos (nodes[558], nodes[211],  nodes[138]);
    nmos (nodes[558], nodes[211],  nodes[138]);
    nmos (nodes[1027], nodes[1649],  nodes[943]);
    nmos (nodes[187], nodes[558],  nodes[926]);
    nmos (nodes[604], nodes[1118],  nodes[638]);
    nmos (nodes[558], nodes[396],  nodes[1358]);
    nmos (nodes[435], nodes[657],  nodes[634]);
    nmos (nodes[435], nodes[657],  nodes[634]);
    nmos (nodes[435], nodes[657],  nodes[634]);
    nmos (nodes[435], nodes[657],  nodes[634]);
    nmos (nodes[657], nodes[435],  nodes[634]);
    nmos (nodes[1568], nodes[1099],  nodes[1542]);
    nmos (nodes[1498], nodes[1184],  nodes[1253]);
    nmos (nodes[558], nodes[903],  nodes[1253]);
    nmos (nodes[1471], nodes[558],  nodes[827]);
    nmos (nodes[558], nodes[392],  nodes[386]);
    nmos (nodes[558], nodes[1704],  nodes[386]);
    nmos (nodes[1565], nodes[700],  nodes[943]);
    nmos (nodes[558], nodes[1166],  nodes[329]);
    nmos (nodes[558], nodes[1704],  nodes[329]);
    nmos (nodes[558], nodes[1107],  nodes[492]);
    nmos (nodes[558], nodes[1005],  nodes[1072]);
    nmos (nodes[1005], nodes[558],  nodes[1072]);
    nmos (nodes[558], nodes[1005],  nodes[1072]);
    nmos (nodes[1005], nodes[558],  nodes[1072]);
    nmos (nodes[558], nodes[1005],  nodes[1072]);
    nmos (nodes[1005], nodes[558],  nodes[1072]);
    nmos (nodes[558], nodes[1005],  nodes[1072]);
    nmos (nodes[1005], nodes[558],  nodes[1072]);
    nmos (nodes[547], nodes[486],  nodes[1571]);
    nmos (nodes[558], nodes[817],  nodes[1571]);
    nmos (nodes[657], nodes[230],  nodes[826]);
    nmos (nodes[1716], nodes[558],  nodes[218]);
    nmos (nodes[688], nodes[1594],  nodes[943]);
    nmos (nodes[67], nodes[558],  nodes[1395]);
    nmos (nodes[558], nodes[67],  nodes[1395]);
    nmos (nodes[1111], nodes[941],  nodes[215]);
    nmos (nodes[250], nodes[155],  nodes[59]);
    nmos (nodes[669], nodes[558],  nodes[1504]);
    nmos (nodes[282], nodes[558],  nodes[6]);
    nmos (nodes[657], nodes[874],  nodes[6]);
    nmos (nodes[1037], nodes[1280],  nodes[145]);
    nmos (nodes[558], nodes[35],  nodes[43]);
    nmos (nodes[583], nodes[558],  nodes[991]);
    nmos (nodes[558], nodes[730],  nodes[448]);
    nmos (nodes[1567], nodes[558],  nodes[678]);
    nmos (nodes[1319], nodes[361],  nodes[943]);
    nmos (nodes[93], nodes[758],  nodes[943]);
    nmos (nodes[558], nodes[1152],  nodes[951]);
    nmos (nodes[657], nodes[642],  nodes[951]);
    nmos (nodes[657], nodes[1287],  nodes[943]);
    nmos (nodes[752], nodes[1190],  nodes[943]);
    nmos (nodes[657], nodes[892],  nodes[943]);
    nmos (nodes[558], nodes[1130],  nodes[1258]);
    nmos (nodes[586], nodes[558],  nodes[1619]);
    nmos (nodes[558], nodes[356],  nodes[923]);
    nmos (nodes[558], nodes[1334],  nodes[923]);
    nmos (nodes[558], nodes[810],  nodes[923]);
    

    supply0 gnd;
    supply1 vcc;
    assign nodes[558] = gnd;
    assign nodes[657] = vcc;

    assign reset  = nodes[159],
           ready  = nodes[89],
           clock0 = nodes[1171],
           clock1 = nodes[1163],
           clock2 = nodes[421],
           irq    = nodes[103], 
           nmi    = nodes[1297],
           so     = nodes[1672];
     //      sync   =  nodes[];

     assign readNotWrite = nodes[1156] ;
     assign address = {
         nodes[195], 
         nodes[672], 
         nodes[349], 
         nodes[1237], 
         nodes[399], 
         nodes[1443], 
         nodes[148], 
         nodes[230], 
         nodes[1493], 
         nodes[887], 
         nodes[736], 
         nodes[435], 
         nodes[211], 
         nodes[1340], 
         nodes[451], 
         nodes[268]
         
     };

     assign data = {
         nodes[1349], 
         nodes[1591], 
         nodes[175], 
         nodes[1393], 
         nodes[650], 
         nodes[945], 
         nodes[82], 
         nodes[1005]
         
     };

endmodule
